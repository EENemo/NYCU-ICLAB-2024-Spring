# 
#              Synchronous High Speed Single Port SRAM Compiler 
# 
#                    UMC 0.18um GenericII Logic Process
#    __________________________________________________________________________
# 
# 
#      (C) Copyright 2002-2009 Faraday Technology Corp. All Rights Reserved.
#    
#    This source code is an unpublished work belongs to Faraday Technology
#    Corp.  It is considered a trade secret and is not to be divulged or
#    used by parties who have not received written authorization from
#    Faraday Technology Corp.
#    
#    Faraday's home page can be found at:
#    http://www.faraday-tech.com/
#   
#       Module Name      : SUMA_400_M1
#       Words            : 400
#       Bits             : 8
#       Byte-Write       : 1
#       Aspect Ratio     : 1
#       Output Loading   : 0.05  (pf)
#       Data Slew        : 0.02  (ns)
#       CK Slew          : 0.02  (ns)
#       Power Ring Width : 2  (um)
# 
# -----------------------------------------------------------------------------
# 
#       Library          : FSA0M_A
#       Memaker          : 200901.2.1
#       Date             : 2024/03/30 23:41:54
# 
# -----------------------------------------------------------------------------


NAMESCASESENSITIVE ON ;
MACRO SUMA_400_M1
CLASS BLOCK ;
FOREIGN SUMA_400_M1 0.000 0.000 ;
ORIGIN 0.000 0.000 ;
SIZE 213.900 BY 259.840 ;
SYMMETRY x y r90 ;
SITE core ;
PIN GND
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
 PORT
  LAYER ME4 ;
  RECT 212.780 247.300 213.900 250.540 ;
  LAYER ME3 ;
  RECT 212.780 247.300 213.900 250.540 ;
  LAYER ME2 ;
  RECT 212.780 247.300 213.900 250.540 ;
  LAYER ME1 ;
  RECT 212.780 247.300 213.900 250.540 ;
 END
 PORT
  LAYER ME4 ;
  RECT 212.780 208.100 213.900 211.340 ;
  LAYER ME3 ;
  RECT 212.780 208.100 213.900 211.340 ;
  LAYER ME2 ;
  RECT 212.780 208.100 213.900 211.340 ;
  LAYER ME1 ;
  RECT 212.780 208.100 213.900 211.340 ;
 END
 PORT
  LAYER ME4 ;
  RECT 212.780 200.260 213.900 203.500 ;
  LAYER ME3 ;
  RECT 212.780 200.260 213.900 203.500 ;
  LAYER ME2 ;
  RECT 212.780 200.260 213.900 203.500 ;
  LAYER ME1 ;
  RECT 212.780 200.260 213.900 203.500 ;
 END
 PORT
  LAYER ME4 ;
  RECT 212.780 192.420 213.900 195.660 ;
  LAYER ME3 ;
  RECT 212.780 192.420 213.900 195.660 ;
  LAYER ME2 ;
  RECT 212.780 192.420 213.900 195.660 ;
  LAYER ME1 ;
  RECT 212.780 192.420 213.900 195.660 ;
 END
 PORT
  LAYER ME4 ;
  RECT 212.780 184.580 213.900 187.820 ;
  LAYER ME3 ;
  RECT 212.780 184.580 213.900 187.820 ;
  LAYER ME2 ;
  RECT 212.780 184.580 213.900 187.820 ;
  LAYER ME1 ;
  RECT 212.780 184.580 213.900 187.820 ;
 END
 PORT
  LAYER ME4 ;
  RECT 212.780 176.740 213.900 179.980 ;
  LAYER ME3 ;
  RECT 212.780 176.740 213.900 179.980 ;
  LAYER ME2 ;
  RECT 212.780 176.740 213.900 179.980 ;
  LAYER ME1 ;
  RECT 212.780 176.740 213.900 179.980 ;
 END
 PORT
  LAYER ME4 ;
  RECT 212.780 168.900 213.900 172.140 ;
  LAYER ME3 ;
  RECT 212.780 168.900 213.900 172.140 ;
  LAYER ME2 ;
  RECT 212.780 168.900 213.900 172.140 ;
  LAYER ME1 ;
  RECT 212.780 168.900 213.900 172.140 ;
 END
 PORT
  LAYER ME4 ;
  RECT 212.780 129.700 213.900 132.940 ;
  LAYER ME3 ;
  RECT 212.780 129.700 213.900 132.940 ;
  LAYER ME2 ;
  RECT 212.780 129.700 213.900 132.940 ;
  LAYER ME1 ;
  RECT 212.780 129.700 213.900 132.940 ;
 END
 PORT
  LAYER ME4 ;
  RECT 212.780 121.860 213.900 125.100 ;
  LAYER ME3 ;
  RECT 212.780 121.860 213.900 125.100 ;
  LAYER ME2 ;
  RECT 212.780 121.860 213.900 125.100 ;
  LAYER ME1 ;
  RECT 212.780 121.860 213.900 125.100 ;
 END
 PORT
  LAYER ME4 ;
  RECT 212.780 114.020 213.900 117.260 ;
  LAYER ME3 ;
  RECT 212.780 114.020 213.900 117.260 ;
  LAYER ME2 ;
  RECT 212.780 114.020 213.900 117.260 ;
  LAYER ME1 ;
  RECT 212.780 114.020 213.900 117.260 ;
 END
 PORT
  LAYER ME4 ;
  RECT 212.780 106.180 213.900 109.420 ;
  LAYER ME3 ;
  RECT 212.780 106.180 213.900 109.420 ;
  LAYER ME2 ;
  RECT 212.780 106.180 213.900 109.420 ;
  LAYER ME1 ;
  RECT 212.780 106.180 213.900 109.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 212.780 98.340 213.900 101.580 ;
  LAYER ME3 ;
  RECT 212.780 98.340 213.900 101.580 ;
  LAYER ME2 ;
  RECT 212.780 98.340 213.900 101.580 ;
  LAYER ME1 ;
  RECT 212.780 98.340 213.900 101.580 ;
 END
 PORT
  LAYER ME4 ;
  RECT 212.780 90.500 213.900 93.740 ;
  LAYER ME3 ;
  RECT 212.780 90.500 213.900 93.740 ;
  LAYER ME2 ;
  RECT 212.780 90.500 213.900 93.740 ;
  LAYER ME1 ;
  RECT 212.780 90.500 213.900 93.740 ;
 END
 PORT
  LAYER ME4 ;
  RECT 212.780 51.300 213.900 54.540 ;
  LAYER ME3 ;
  RECT 212.780 51.300 213.900 54.540 ;
  LAYER ME2 ;
  RECT 212.780 51.300 213.900 54.540 ;
  LAYER ME1 ;
  RECT 212.780 51.300 213.900 54.540 ;
 END
 PORT
  LAYER ME4 ;
  RECT 212.780 43.460 213.900 46.700 ;
  LAYER ME3 ;
  RECT 212.780 43.460 213.900 46.700 ;
  LAYER ME2 ;
  RECT 212.780 43.460 213.900 46.700 ;
  LAYER ME1 ;
  RECT 212.780 43.460 213.900 46.700 ;
 END
 PORT
  LAYER ME4 ;
  RECT 212.780 35.620 213.900 38.860 ;
  LAYER ME3 ;
  RECT 212.780 35.620 213.900 38.860 ;
  LAYER ME2 ;
  RECT 212.780 35.620 213.900 38.860 ;
  LAYER ME1 ;
  RECT 212.780 35.620 213.900 38.860 ;
 END
 PORT
  LAYER ME4 ;
  RECT 212.780 27.780 213.900 31.020 ;
  LAYER ME3 ;
  RECT 212.780 27.780 213.900 31.020 ;
  LAYER ME2 ;
  RECT 212.780 27.780 213.900 31.020 ;
  LAYER ME1 ;
  RECT 212.780 27.780 213.900 31.020 ;
 END
 PORT
  LAYER ME4 ;
  RECT 212.780 19.940 213.900 23.180 ;
  LAYER ME3 ;
  RECT 212.780 19.940 213.900 23.180 ;
  LAYER ME2 ;
  RECT 212.780 19.940 213.900 23.180 ;
  LAYER ME1 ;
  RECT 212.780 19.940 213.900 23.180 ;
 END
 PORT
  LAYER ME4 ;
  RECT 212.780 12.100 213.900 15.340 ;
  LAYER ME3 ;
  RECT 212.780 12.100 213.900 15.340 ;
  LAYER ME2 ;
  RECT 212.780 12.100 213.900 15.340 ;
  LAYER ME1 ;
  RECT 212.780 12.100 213.900 15.340 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 247.300 1.120 250.540 ;
  LAYER ME3 ;
  RECT 0.000 247.300 1.120 250.540 ;
  LAYER ME2 ;
  RECT 0.000 247.300 1.120 250.540 ;
  LAYER ME1 ;
  RECT 0.000 247.300 1.120 250.540 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 208.100 1.120 211.340 ;
  LAYER ME3 ;
  RECT 0.000 208.100 1.120 211.340 ;
  LAYER ME2 ;
  RECT 0.000 208.100 1.120 211.340 ;
  LAYER ME1 ;
  RECT 0.000 208.100 1.120 211.340 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 200.260 1.120 203.500 ;
  LAYER ME3 ;
  RECT 0.000 200.260 1.120 203.500 ;
  LAYER ME2 ;
  RECT 0.000 200.260 1.120 203.500 ;
  LAYER ME1 ;
  RECT 0.000 200.260 1.120 203.500 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 192.420 1.120 195.660 ;
  LAYER ME3 ;
  RECT 0.000 192.420 1.120 195.660 ;
  LAYER ME2 ;
  RECT 0.000 192.420 1.120 195.660 ;
  LAYER ME1 ;
  RECT 0.000 192.420 1.120 195.660 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 184.580 1.120 187.820 ;
  LAYER ME3 ;
  RECT 0.000 184.580 1.120 187.820 ;
  LAYER ME2 ;
  RECT 0.000 184.580 1.120 187.820 ;
  LAYER ME1 ;
  RECT 0.000 184.580 1.120 187.820 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 176.740 1.120 179.980 ;
  LAYER ME3 ;
  RECT 0.000 176.740 1.120 179.980 ;
  LAYER ME2 ;
  RECT 0.000 176.740 1.120 179.980 ;
  LAYER ME1 ;
  RECT 0.000 176.740 1.120 179.980 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 168.900 1.120 172.140 ;
  LAYER ME3 ;
  RECT 0.000 168.900 1.120 172.140 ;
  LAYER ME2 ;
  RECT 0.000 168.900 1.120 172.140 ;
  LAYER ME1 ;
  RECT 0.000 168.900 1.120 172.140 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 129.700 1.120 132.940 ;
  LAYER ME3 ;
  RECT 0.000 129.700 1.120 132.940 ;
  LAYER ME2 ;
  RECT 0.000 129.700 1.120 132.940 ;
  LAYER ME1 ;
  RECT 0.000 129.700 1.120 132.940 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 121.860 1.120 125.100 ;
  LAYER ME3 ;
  RECT 0.000 121.860 1.120 125.100 ;
  LAYER ME2 ;
  RECT 0.000 121.860 1.120 125.100 ;
  LAYER ME1 ;
  RECT 0.000 121.860 1.120 125.100 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 114.020 1.120 117.260 ;
  LAYER ME3 ;
  RECT 0.000 114.020 1.120 117.260 ;
  LAYER ME2 ;
  RECT 0.000 114.020 1.120 117.260 ;
  LAYER ME1 ;
  RECT 0.000 114.020 1.120 117.260 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 106.180 1.120 109.420 ;
  LAYER ME3 ;
  RECT 0.000 106.180 1.120 109.420 ;
  LAYER ME2 ;
  RECT 0.000 106.180 1.120 109.420 ;
  LAYER ME1 ;
  RECT 0.000 106.180 1.120 109.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 98.340 1.120 101.580 ;
  LAYER ME3 ;
  RECT 0.000 98.340 1.120 101.580 ;
  LAYER ME2 ;
  RECT 0.000 98.340 1.120 101.580 ;
  LAYER ME1 ;
  RECT 0.000 98.340 1.120 101.580 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 90.500 1.120 93.740 ;
  LAYER ME3 ;
  RECT 0.000 90.500 1.120 93.740 ;
  LAYER ME2 ;
  RECT 0.000 90.500 1.120 93.740 ;
  LAYER ME1 ;
  RECT 0.000 90.500 1.120 93.740 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 51.300 1.120 54.540 ;
  LAYER ME3 ;
  RECT 0.000 51.300 1.120 54.540 ;
  LAYER ME2 ;
  RECT 0.000 51.300 1.120 54.540 ;
  LAYER ME1 ;
  RECT 0.000 51.300 1.120 54.540 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 43.460 1.120 46.700 ;
  LAYER ME3 ;
  RECT 0.000 43.460 1.120 46.700 ;
  LAYER ME2 ;
  RECT 0.000 43.460 1.120 46.700 ;
  LAYER ME1 ;
  RECT 0.000 43.460 1.120 46.700 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 35.620 1.120 38.860 ;
  LAYER ME3 ;
  RECT 0.000 35.620 1.120 38.860 ;
  LAYER ME2 ;
  RECT 0.000 35.620 1.120 38.860 ;
  LAYER ME1 ;
  RECT 0.000 35.620 1.120 38.860 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 27.780 1.120 31.020 ;
  LAYER ME3 ;
  RECT 0.000 27.780 1.120 31.020 ;
  LAYER ME2 ;
  RECT 0.000 27.780 1.120 31.020 ;
  LAYER ME1 ;
  RECT 0.000 27.780 1.120 31.020 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 19.940 1.120 23.180 ;
  LAYER ME3 ;
  RECT 0.000 19.940 1.120 23.180 ;
  LAYER ME2 ;
  RECT 0.000 19.940 1.120 23.180 ;
  LAYER ME1 ;
  RECT 0.000 19.940 1.120 23.180 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 12.100 1.120 15.340 ;
  LAYER ME3 ;
  RECT 0.000 12.100 1.120 15.340 ;
  LAYER ME2 ;
  RECT 0.000 12.100 1.120 15.340 ;
  LAYER ME1 ;
  RECT 0.000 12.100 1.120 15.340 ;
 END
 PORT
  LAYER ME4 ;
  RECT 194.460 258.720 198.000 259.840 ;
  LAYER ME3 ;
  RECT 194.460 258.720 198.000 259.840 ;
  LAYER ME2 ;
  RECT 194.460 258.720 198.000 259.840 ;
  LAYER ME1 ;
  RECT 194.460 258.720 198.000 259.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 185.780 258.720 189.320 259.840 ;
  LAYER ME3 ;
  RECT 185.780 258.720 189.320 259.840 ;
  LAYER ME2 ;
  RECT 185.780 258.720 189.320 259.840 ;
  LAYER ME1 ;
  RECT 185.780 258.720 189.320 259.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 142.380 258.720 145.920 259.840 ;
  LAYER ME3 ;
  RECT 142.380 258.720 145.920 259.840 ;
  LAYER ME2 ;
  RECT 142.380 258.720 145.920 259.840 ;
  LAYER ME1 ;
  RECT 142.380 258.720 145.920 259.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 133.700 258.720 137.240 259.840 ;
  LAYER ME3 ;
  RECT 133.700 258.720 137.240 259.840 ;
  LAYER ME2 ;
  RECT 133.700 258.720 137.240 259.840 ;
  LAYER ME1 ;
  RECT 133.700 258.720 137.240 259.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 125.020 258.720 128.560 259.840 ;
  LAYER ME3 ;
  RECT 125.020 258.720 128.560 259.840 ;
  LAYER ME2 ;
  RECT 125.020 258.720 128.560 259.840 ;
  LAYER ME1 ;
  RECT 125.020 258.720 128.560 259.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 116.340 258.720 119.880 259.840 ;
  LAYER ME3 ;
  RECT 116.340 258.720 119.880 259.840 ;
  LAYER ME2 ;
  RECT 116.340 258.720 119.880 259.840 ;
  LAYER ME1 ;
  RECT 116.340 258.720 119.880 259.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 107.660 258.720 111.200 259.840 ;
  LAYER ME3 ;
  RECT 107.660 258.720 111.200 259.840 ;
  LAYER ME2 ;
  RECT 107.660 258.720 111.200 259.840 ;
  LAYER ME1 ;
  RECT 107.660 258.720 111.200 259.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 98.980 258.720 102.520 259.840 ;
  LAYER ME3 ;
  RECT 98.980 258.720 102.520 259.840 ;
  LAYER ME2 ;
  RECT 98.980 258.720 102.520 259.840 ;
  LAYER ME1 ;
  RECT 98.980 258.720 102.520 259.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 55.580 258.720 59.120 259.840 ;
  LAYER ME3 ;
  RECT 55.580 258.720 59.120 259.840 ;
  LAYER ME2 ;
  RECT 55.580 258.720 59.120 259.840 ;
  LAYER ME1 ;
  RECT 55.580 258.720 59.120 259.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 46.900 258.720 50.440 259.840 ;
  LAYER ME3 ;
  RECT 46.900 258.720 50.440 259.840 ;
  LAYER ME2 ;
  RECT 46.900 258.720 50.440 259.840 ;
  LAYER ME1 ;
  RECT 46.900 258.720 50.440 259.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 38.220 258.720 41.760 259.840 ;
  LAYER ME3 ;
  RECT 38.220 258.720 41.760 259.840 ;
  LAYER ME2 ;
  RECT 38.220 258.720 41.760 259.840 ;
  LAYER ME1 ;
  RECT 38.220 258.720 41.760 259.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 29.540 258.720 33.080 259.840 ;
  LAYER ME3 ;
  RECT 29.540 258.720 33.080 259.840 ;
  LAYER ME2 ;
  RECT 29.540 258.720 33.080 259.840 ;
  LAYER ME1 ;
  RECT 29.540 258.720 33.080 259.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 20.860 258.720 24.400 259.840 ;
  LAYER ME3 ;
  RECT 20.860 258.720 24.400 259.840 ;
  LAYER ME2 ;
  RECT 20.860 258.720 24.400 259.840 ;
  LAYER ME1 ;
  RECT 20.860 258.720 24.400 259.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 12.180 258.720 15.720 259.840 ;
  LAYER ME3 ;
  RECT 12.180 258.720 15.720 259.840 ;
  LAYER ME2 ;
  RECT 12.180 258.720 15.720 259.840 ;
  LAYER ME1 ;
  RECT 12.180 258.720 15.720 259.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 119.440 0.000 122.980 1.120 ;
  LAYER ME3 ;
  RECT 119.440 0.000 122.980 1.120 ;
  LAYER ME2 ;
  RECT 119.440 0.000 122.980 1.120 ;
  LAYER ME1 ;
  RECT 119.440 0.000 122.980 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 97.740 0.000 101.280 1.120 ;
  LAYER ME3 ;
  RECT 97.740 0.000 101.280 1.120 ;
  LAYER ME2 ;
  RECT 97.740 0.000 101.280 1.120 ;
  LAYER ME1 ;
  RECT 97.740 0.000 101.280 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 76.660 0.000 80.200 1.120 ;
  LAYER ME3 ;
  RECT 76.660 0.000 80.200 1.120 ;
  LAYER ME2 ;
  RECT 76.660 0.000 80.200 1.120 ;
  LAYER ME1 ;
  RECT 76.660 0.000 80.200 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 65.500 0.000 69.040 1.120 ;
  LAYER ME3 ;
  RECT 65.500 0.000 69.040 1.120 ;
  LAYER ME2 ;
  RECT 65.500 0.000 69.040 1.120 ;
  LAYER ME1 ;
  RECT 65.500 0.000 69.040 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 43.800 0.000 47.340 1.120 ;
  LAYER ME3 ;
  RECT 43.800 0.000 47.340 1.120 ;
  LAYER ME2 ;
  RECT 43.800 0.000 47.340 1.120 ;
  LAYER ME1 ;
  RECT 43.800 0.000 47.340 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 27.060 0.000 30.600 1.120 ;
  LAYER ME3 ;
  RECT 27.060 0.000 30.600 1.120 ;
  LAYER ME2 ;
  RECT 27.060 0.000 30.600 1.120 ;
  LAYER ME1 ;
  RECT 27.060 0.000 30.600 1.120 ;
 END
END GND
PIN VCC
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
 PORT
  LAYER ME4 ;
  RECT 212.780 243.380 213.900 246.620 ;
  LAYER ME3 ;
  RECT 212.780 243.380 213.900 246.620 ;
  LAYER ME2 ;
  RECT 212.780 243.380 213.900 246.620 ;
  LAYER ME1 ;
  RECT 212.780 243.380 213.900 246.620 ;
 END
 PORT
  LAYER ME4 ;
  RECT 212.780 204.180 213.900 207.420 ;
  LAYER ME3 ;
  RECT 212.780 204.180 213.900 207.420 ;
  LAYER ME2 ;
  RECT 212.780 204.180 213.900 207.420 ;
  LAYER ME1 ;
  RECT 212.780 204.180 213.900 207.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 212.780 196.340 213.900 199.580 ;
  LAYER ME3 ;
  RECT 212.780 196.340 213.900 199.580 ;
  LAYER ME2 ;
  RECT 212.780 196.340 213.900 199.580 ;
  LAYER ME1 ;
  RECT 212.780 196.340 213.900 199.580 ;
 END
 PORT
  LAYER ME4 ;
  RECT 212.780 188.500 213.900 191.740 ;
  LAYER ME3 ;
  RECT 212.780 188.500 213.900 191.740 ;
  LAYER ME2 ;
  RECT 212.780 188.500 213.900 191.740 ;
  LAYER ME1 ;
  RECT 212.780 188.500 213.900 191.740 ;
 END
 PORT
  LAYER ME4 ;
  RECT 212.780 180.660 213.900 183.900 ;
  LAYER ME3 ;
  RECT 212.780 180.660 213.900 183.900 ;
  LAYER ME2 ;
  RECT 212.780 180.660 213.900 183.900 ;
  LAYER ME1 ;
  RECT 212.780 180.660 213.900 183.900 ;
 END
 PORT
  LAYER ME4 ;
  RECT 212.780 172.820 213.900 176.060 ;
  LAYER ME3 ;
  RECT 212.780 172.820 213.900 176.060 ;
  LAYER ME2 ;
  RECT 212.780 172.820 213.900 176.060 ;
  LAYER ME1 ;
  RECT 212.780 172.820 213.900 176.060 ;
 END
 PORT
  LAYER ME4 ;
  RECT 212.780 164.980 213.900 168.220 ;
  LAYER ME3 ;
  RECT 212.780 164.980 213.900 168.220 ;
  LAYER ME2 ;
  RECT 212.780 164.980 213.900 168.220 ;
  LAYER ME1 ;
  RECT 212.780 164.980 213.900 168.220 ;
 END
 PORT
  LAYER ME4 ;
  RECT 212.780 125.780 213.900 129.020 ;
  LAYER ME3 ;
  RECT 212.780 125.780 213.900 129.020 ;
  LAYER ME2 ;
  RECT 212.780 125.780 213.900 129.020 ;
  LAYER ME1 ;
  RECT 212.780 125.780 213.900 129.020 ;
 END
 PORT
  LAYER ME4 ;
  RECT 212.780 117.940 213.900 121.180 ;
  LAYER ME3 ;
  RECT 212.780 117.940 213.900 121.180 ;
  LAYER ME2 ;
  RECT 212.780 117.940 213.900 121.180 ;
  LAYER ME1 ;
  RECT 212.780 117.940 213.900 121.180 ;
 END
 PORT
  LAYER ME4 ;
  RECT 212.780 110.100 213.900 113.340 ;
  LAYER ME3 ;
  RECT 212.780 110.100 213.900 113.340 ;
  LAYER ME2 ;
  RECT 212.780 110.100 213.900 113.340 ;
  LAYER ME1 ;
  RECT 212.780 110.100 213.900 113.340 ;
 END
 PORT
  LAYER ME4 ;
  RECT 212.780 102.260 213.900 105.500 ;
  LAYER ME3 ;
  RECT 212.780 102.260 213.900 105.500 ;
  LAYER ME2 ;
  RECT 212.780 102.260 213.900 105.500 ;
  LAYER ME1 ;
  RECT 212.780 102.260 213.900 105.500 ;
 END
 PORT
  LAYER ME4 ;
  RECT 212.780 94.420 213.900 97.660 ;
  LAYER ME3 ;
  RECT 212.780 94.420 213.900 97.660 ;
  LAYER ME2 ;
  RECT 212.780 94.420 213.900 97.660 ;
  LAYER ME1 ;
  RECT 212.780 94.420 213.900 97.660 ;
 END
 PORT
  LAYER ME4 ;
  RECT 212.780 86.580 213.900 89.820 ;
  LAYER ME3 ;
  RECT 212.780 86.580 213.900 89.820 ;
  LAYER ME2 ;
  RECT 212.780 86.580 213.900 89.820 ;
  LAYER ME1 ;
  RECT 212.780 86.580 213.900 89.820 ;
 END
 PORT
  LAYER ME4 ;
  RECT 212.780 47.380 213.900 50.620 ;
  LAYER ME3 ;
  RECT 212.780 47.380 213.900 50.620 ;
  LAYER ME2 ;
  RECT 212.780 47.380 213.900 50.620 ;
  LAYER ME1 ;
  RECT 212.780 47.380 213.900 50.620 ;
 END
 PORT
  LAYER ME4 ;
  RECT 212.780 39.540 213.900 42.780 ;
  LAYER ME3 ;
  RECT 212.780 39.540 213.900 42.780 ;
  LAYER ME2 ;
  RECT 212.780 39.540 213.900 42.780 ;
  LAYER ME1 ;
  RECT 212.780 39.540 213.900 42.780 ;
 END
 PORT
  LAYER ME4 ;
  RECT 212.780 31.700 213.900 34.940 ;
  LAYER ME3 ;
  RECT 212.780 31.700 213.900 34.940 ;
  LAYER ME2 ;
  RECT 212.780 31.700 213.900 34.940 ;
  LAYER ME1 ;
  RECT 212.780 31.700 213.900 34.940 ;
 END
 PORT
  LAYER ME4 ;
  RECT 212.780 23.860 213.900 27.100 ;
  LAYER ME3 ;
  RECT 212.780 23.860 213.900 27.100 ;
  LAYER ME2 ;
  RECT 212.780 23.860 213.900 27.100 ;
  LAYER ME1 ;
  RECT 212.780 23.860 213.900 27.100 ;
 END
 PORT
  LAYER ME4 ;
  RECT 212.780 16.020 213.900 19.260 ;
  LAYER ME3 ;
  RECT 212.780 16.020 213.900 19.260 ;
  LAYER ME2 ;
  RECT 212.780 16.020 213.900 19.260 ;
  LAYER ME1 ;
  RECT 212.780 16.020 213.900 19.260 ;
 END
 PORT
  LAYER ME4 ;
  RECT 212.780 8.180 213.900 11.420 ;
  LAYER ME3 ;
  RECT 212.780 8.180 213.900 11.420 ;
  LAYER ME2 ;
  RECT 212.780 8.180 213.900 11.420 ;
  LAYER ME1 ;
  RECT 212.780 8.180 213.900 11.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 243.380 1.120 246.620 ;
  LAYER ME3 ;
  RECT 0.000 243.380 1.120 246.620 ;
  LAYER ME2 ;
  RECT 0.000 243.380 1.120 246.620 ;
  LAYER ME1 ;
  RECT 0.000 243.380 1.120 246.620 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 204.180 1.120 207.420 ;
  LAYER ME3 ;
  RECT 0.000 204.180 1.120 207.420 ;
  LAYER ME2 ;
  RECT 0.000 204.180 1.120 207.420 ;
  LAYER ME1 ;
  RECT 0.000 204.180 1.120 207.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 196.340 1.120 199.580 ;
  LAYER ME3 ;
  RECT 0.000 196.340 1.120 199.580 ;
  LAYER ME2 ;
  RECT 0.000 196.340 1.120 199.580 ;
  LAYER ME1 ;
  RECT 0.000 196.340 1.120 199.580 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 188.500 1.120 191.740 ;
  LAYER ME3 ;
  RECT 0.000 188.500 1.120 191.740 ;
  LAYER ME2 ;
  RECT 0.000 188.500 1.120 191.740 ;
  LAYER ME1 ;
  RECT 0.000 188.500 1.120 191.740 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 180.660 1.120 183.900 ;
  LAYER ME3 ;
  RECT 0.000 180.660 1.120 183.900 ;
  LAYER ME2 ;
  RECT 0.000 180.660 1.120 183.900 ;
  LAYER ME1 ;
  RECT 0.000 180.660 1.120 183.900 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 172.820 1.120 176.060 ;
  LAYER ME3 ;
  RECT 0.000 172.820 1.120 176.060 ;
  LAYER ME2 ;
  RECT 0.000 172.820 1.120 176.060 ;
  LAYER ME1 ;
  RECT 0.000 172.820 1.120 176.060 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 164.980 1.120 168.220 ;
  LAYER ME3 ;
  RECT 0.000 164.980 1.120 168.220 ;
  LAYER ME2 ;
  RECT 0.000 164.980 1.120 168.220 ;
  LAYER ME1 ;
  RECT 0.000 164.980 1.120 168.220 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 125.780 1.120 129.020 ;
  LAYER ME3 ;
  RECT 0.000 125.780 1.120 129.020 ;
  LAYER ME2 ;
  RECT 0.000 125.780 1.120 129.020 ;
  LAYER ME1 ;
  RECT 0.000 125.780 1.120 129.020 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 117.940 1.120 121.180 ;
  LAYER ME3 ;
  RECT 0.000 117.940 1.120 121.180 ;
  LAYER ME2 ;
  RECT 0.000 117.940 1.120 121.180 ;
  LAYER ME1 ;
  RECT 0.000 117.940 1.120 121.180 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 110.100 1.120 113.340 ;
  LAYER ME3 ;
  RECT 0.000 110.100 1.120 113.340 ;
  LAYER ME2 ;
  RECT 0.000 110.100 1.120 113.340 ;
  LAYER ME1 ;
  RECT 0.000 110.100 1.120 113.340 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 102.260 1.120 105.500 ;
  LAYER ME3 ;
  RECT 0.000 102.260 1.120 105.500 ;
  LAYER ME2 ;
  RECT 0.000 102.260 1.120 105.500 ;
  LAYER ME1 ;
  RECT 0.000 102.260 1.120 105.500 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 94.420 1.120 97.660 ;
  LAYER ME3 ;
  RECT 0.000 94.420 1.120 97.660 ;
  LAYER ME2 ;
  RECT 0.000 94.420 1.120 97.660 ;
  LAYER ME1 ;
  RECT 0.000 94.420 1.120 97.660 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 86.580 1.120 89.820 ;
  LAYER ME3 ;
  RECT 0.000 86.580 1.120 89.820 ;
  LAYER ME2 ;
  RECT 0.000 86.580 1.120 89.820 ;
  LAYER ME1 ;
  RECT 0.000 86.580 1.120 89.820 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 47.380 1.120 50.620 ;
  LAYER ME3 ;
  RECT 0.000 47.380 1.120 50.620 ;
  LAYER ME2 ;
  RECT 0.000 47.380 1.120 50.620 ;
  LAYER ME1 ;
  RECT 0.000 47.380 1.120 50.620 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 39.540 1.120 42.780 ;
  LAYER ME3 ;
  RECT 0.000 39.540 1.120 42.780 ;
  LAYER ME2 ;
  RECT 0.000 39.540 1.120 42.780 ;
  LAYER ME1 ;
  RECT 0.000 39.540 1.120 42.780 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 31.700 1.120 34.940 ;
  LAYER ME3 ;
  RECT 0.000 31.700 1.120 34.940 ;
  LAYER ME2 ;
  RECT 0.000 31.700 1.120 34.940 ;
  LAYER ME1 ;
  RECT 0.000 31.700 1.120 34.940 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 23.860 1.120 27.100 ;
  LAYER ME3 ;
  RECT 0.000 23.860 1.120 27.100 ;
  LAYER ME2 ;
  RECT 0.000 23.860 1.120 27.100 ;
  LAYER ME1 ;
  RECT 0.000 23.860 1.120 27.100 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 16.020 1.120 19.260 ;
  LAYER ME3 ;
  RECT 0.000 16.020 1.120 19.260 ;
  LAYER ME2 ;
  RECT 0.000 16.020 1.120 19.260 ;
  LAYER ME1 ;
  RECT 0.000 16.020 1.120 19.260 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 8.180 1.120 11.420 ;
  LAYER ME3 ;
  RECT 0.000 8.180 1.120 11.420 ;
  LAYER ME2 ;
  RECT 0.000 8.180 1.120 11.420 ;
  LAYER ME1 ;
  RECT 0.000 8.180 1.120 11.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 198.800 258.720 202.340 259.840 ;
  LAYER ME3 ;
  RECT 198.800 258.720 202.340 259.840 ;
  LAYER ME2 ;
  RECT 198.800 258.720 202.340 259.840 ;
  LAYER ME1 ;
  RECT 198.800 258.720 202.340 259.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 190.120 258.720 193.660 259.840 ;
  LAYER ME3 ;
  RECT 190.120 258.720 193.660 259.840 ;
  LAYER ME2 ;
  RECT 190.120 258.720 193.660 259.840 ;
  LAYER ME1 ;
  RECT 190.120 258.720 193.660 259.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 181.440 258.720 184.980 259.840 ;
  LAYER ME3 ;
  RECT 181.440 258.720 184.980 259.840 ;
  LAYER ME2 ;
  RECT 181.440 258.720 184.980 259.840 ;
  LAYER ME1 ;
  RECT 181.440 258.720 184.980 259.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 138.040 258.720 141.580 259.840 ;
  LAYER ME3 ;
  RECT 138.040 258.720 141.580 259.840 ;
  LAYER ME2 ;
  RECT 138.040 258.720 141.580 259.840 ;
  LAYER ME1 ;
  RECT 138.040 258.720 141.580 259.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 129.360 258.720 132.900 259.840 ;
  LAYER ME3 ;
  RECT 129.360 258.720 132.900 259.840 ;
  LAYER ME2 ;
  RECT 129.360 258.720 132.900 259.840 ;
  LAYER ME1 ;
  RECT 129.360 258.720 132.900 259.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 120.680 258.720 124.220 259.840 ;
  LAYER ME3 ;
  RECT 120.680 258.720 124.220 259.840 ;
  LAYER ME2 ;
  RECT 120.680 258.720 124.220 259.840 ;
  LAYER ME1 ;
  RECT 120.680 258.720 124.220 259.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 112.000 258.720 115.540 259.840 ;
  LAYER ME3 ;
  RECT 112.000 258.720 115.540 259.840 ;
  LAYER ME2 ;
  RECT 112.000 258.720 115.540 259.840 ;
  LAYER ME1 ;
  RECT 112.000 258.720 115.540 259.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 103.320 258.720 106.860 259.840 ;
  LAYER ME3 ;
  RECT 103.320 258.720 106.860 259.840 ;
  LAYER ME2 ;
  RECT 103.320 258.720 106.860 259.840 ;
  LAYER ME1 ;
  RECT 103.320 258.720 106.860 259.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 94.640 258.720 98.180 259.840 ;
  LAYER ME3 ;
  RECT 94.640 258.720 98.180 259.840 ;
  LAYER ME2 ;
  RECT 94.640 258.720 98.180 259.840 ;
  LAYER ME1 ;
  RECT 94.640 258.720 98.180 259.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 51.240 258.720 54.780 259.840 ;
  LAYER ME3 ;
  RECT 51.240 258.720 54.780 259.840 ;
  LAYER ME2 ;
  RECT 51.240 258.720 54.780 259.840 ;
  LAYER ME1 ;
  RECT 51.240 258.720 54.780 259.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 42.560 258.720 46.100 259.840 ;
  LAYER ME3 ;
  RECT 42.560 258.720 46.100 259.840 ;
  LAYER ME2 ;
  RECT 42.560 258.720 46.100 259.840 ;
  LAYER ME1 ;
  RECT 42.560 258.720 46.100 259.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 33.880 258.720 37.420 259.840 ;
  LAYER ME3 ;
  RECT 33.880 258.720 37.420 259.840 ;
  LAYER ME2 ;
  RECT 33.880 258.720 37.420 259.840 ;
  LAYER ME1 ;
  RECT 33.880 258.720 37.420 259.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 25.200 258.720 28.740 259.840 ;
  LAYER ME3 ;
  RECT 25.200 258.720 28.740 259.840 ;
  LAYER ME2 ;
  RECT 25.200 258.720 28.740 259.840 ;
  LAYER ME1 ;
  RECT 25.200 258.720 28.740 259.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 16.520 258.720 20.060 259.840 ;
  LAYER ME3 ;
  RECT 16.520 258.720 20.060 259.840 ;
  LAYER ME2 ;
  RECT 16.520 258.720 20.060 259.840 ;
  LAYER ME1 ;
  RECT 16.520 258.720 20.060 259.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 7.840 258.720 11.380 259.840 ;
  LAYER ME3 ;
  RECT 7.840 258.720 11.380 259.840 ;
  LAYER ME2 ;
  RECT 7.840 258.720 11.380 259.840 ;
  LAYER ME1 ;
  RECT 7.840 258.720 11.380 259.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 115.100 0.000 118.640 1.120 ;
  LAYER ME3 ;
  RECT 115.100 0.000 118.640 1.120 ;
  LAYER ME2 ;
  RECT 115.100 0.000 118.640 1.120 ;
  LAYER ME1 ;
  RECT 115.100 0.000 118.640 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 87.200 0.000 90.740 1.120 ;
  LAYER ME3 ;
  RECT 87.200 0.000 90.740 1.120 ;
  LAYER ME2 ;
  RECT 87.200 0.000 90.740 1.120 ;
  LAYER ME1 ;
  RECT 87.200 0.000 90.740 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 69.840 0.000 73.380 1.120 ;
  LAYER ME3 ;
  RECT 69.840 0.000 73.380 1.120 ;
  LAYER ME2 ;
  RECT 69.840 0.000 73.380 1.120 ;
  LAYER ME1 ;
  RECT 69.840 0.000 73.380 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 56.820 0.000 60.360 1.120 ;
  LAYER ME3 ;
  RECT 56.820 0.000 60.360 1.120 ;
  LAYER ME2 ;
  RECT 56.820 0.000 60.360 1.120 ;
  LAYER ME1 ;
  RECT 56.820 0.000 60.360 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 35.740 0.000 39.280 1.120 ;
  LAYER ME3 ;
  RECT 35.740 0.000 39.280 1.120 ;
  LAYER ME2 ;
  RECT 35.740 0.000 39.280 1.120 ;
  LAYER ME1 ;
  RECT 35.740 0.000 39.280 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 14.040 0.000 17.580 1.120 ;
  LAYER ME3 ;
  RECT 14.040 0.000 17.580 1.120 ;
  LAYER ME2 ;
  RECT 14.040 0.000 17.580 1.120 ;
  LAYER ME1 ;
  RECT 14.040 0.000 17.580 1.120 ;
 END
END VCC
PIN DO7
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 200.320 0.000 201.440 1.120 ;
  LAYER ME3 ;
  RECT 200.320 0.000 201.440 1.120 ;
  LAYER ME2 ;
  RECT 200.320 0.000 201.440 1.120 ;
  LAYER ME1 ;
  RECT 200.320 0.000 201.440 1.120 ;
 END
END DO7
PIN DI7
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 191.640 0.000 192.760 1.120 ;
  LAYER ME3 ;
  RECT 191.640 0.000 192.760 1.120 ;
  LAYER ME2 ;
  RECT 191.640 0.000 192.760 1.120 ;
  LAYER ME1 ;
  RECT 191.640 0.000 192.760 1.120 ;
 END
END DI7
PIN DO6
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 187.300 0.000 188.420 1.120 ;
  LAYER ME3 ;
  RECT 187.300 0.000 188.420 1.120 ;
  LAYER ME2 ;
  RECT 187.300 0.000 188.420 1.120 ;
  LAYER ME1 ;
  RECT 187.300 0.000 188.420 1.120 ;
 END
END DO6
PIN DI6
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 178.620 0.000 179.740 1.120 ;
  LAYER ME3 ;
  RECT 178.620 0.000 179.740 1.120 ;
  LAYER ME2 ;
  RECT 178.620 0.000 179.740 1.120 ;
  LAYER ME1 ;
  RECT 178.620 0.000 179.740 1.120 ;
 END
END DI6
PIN DO5
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 170.560 0.000 171.680 1.120 ;
  LAYER ME3 ;
  RECT 170.560 0.000 171.680 1.120 ;
  LAYER ME2 ;
  RECT 170.560 0.000 171.680 1.120 ;
  LAYER ME1 ;
  RECT 170.560 0.000 171.680 1.120 ;
 END
END DO5
PIN DI5
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 161.880 0.000 163.000 1.120 ;
  LAYER ME3 ;
  RECT 161.880 0.000 163.000 1.120 ;
  LAYER ME2 ;
  RECT 161.880 0.000 163.000 1.120 ;
  LAYER ME1 ;
  RECT 161.880 0.000 163.000 1.120 ;
 END
END DI5
PIN DO4
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 156.920 0.000 158.040 1.120 ;
  LAYER ME3 ;
  RECT 156.920 0.000 158.040 1.120 ;
  LAYER ME2 ;
  RECT 156.920 0.000 158.040 1.120 ;
  LAYER ME1 ;
  RECT 156.920 0.000 158.040 1.120 ;
 END
END DO4
PIN DI4
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 148.860 0.000 149.980 1.120 ;
  LAYER ME3 ;
  RECT 148.860 0.000 149.980 1.120 ;
  LAYER ME2 ;
  RECT 148.860 0.000 149.980 1.120 ;
  LAYER ME1 ;
  RECT 148.860 0.000 149.980 1.120 ;
 END
END DI4
PIN A1
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 143.280 0.000 144.400 1.120 ;
  LAYER ME3 ;
  RECT 143.280 0.000 144.400 1.120 ;
  LAYER ME2 ;
  RECT 143.280 0.000 144.400 1.120 ;
  LAYER ME1 ;
  RECT 143.280 0.000 144.400 1.120 ;
 END
END A1
PIN WEB
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER ME4 ;
  RECT 141.420 0.000 142.540 1.120 ;
  LAYER ME3 ;
  RECT 141.420 0.000 142.540 1.120 ;
  LAYER ME2 ;
  RECT 141.420 0.000 142.540 1.120 ;
  LAYER ME1 ;
  RECT 141.420 0.000 142.540 1.120 ;
 END
END WEB
PIN OE
  DIRECTION INPUT ;
  CAPACITANCE 0.033 ;
 PORT
  LAYER ME4 ;
  RECT 136.460 0.000 137.580 1.120 ;
  LAYER ME3 ;
  RECT 136.460 0.000 137.580 1.120 ;
  LAYER ME2 ;
  RECT 136.460 0.000 137.580 1.120 ;
  LAYER ME1 ;
  RECT 136.460 0.000 137.580 1.120 ;
 END
END OE
PIN CS
  DIRECTION INPUT ;
  CAPACITANCE 0.123 ;
 PORT
  LAYER ME4 ;
  RECT 134.600 0.000 135.720 1.120 ;
  LAYER ME3 ;
  RECT 134.600 0.000 135.720 1.120 ;
  LAYER ME2 ;
  RECT 134.600 0.000 135.720 1.120 ;
  LAYER ME1 ;
  RECT 134.600 0.000 135.720 1.120 ;
 END
END CS
PIN A2
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 112.900 0.000 114.020 1.120 ;
  LAYER ME3 ;
  RECT 112.900 0.000 114.020 1.120 ;
  LAYER ME2 ;
  RECT 112.900 0.000 114.020 1.120 ;
  LAYER ME1 ;
  RECT 112.900 0.000 114.020 1.120 ;
 END
END A2
PIN CK
  DIRECTION INPUT ;
  CAPACITANCE 0.063 ;
 PORT
  LAYER ME4 ;
  RECT 109.800 0.000 110.920 1.120 ;
  LAYER ME3 ;
  RECT 109.800 0.000 110.920 1.120 ;
  LAYER ME2 ;
  RECT 109.800 0.000 110.920 1.120 ;
  LAYER ME1 ;
  RECT 109.800 0.000 110.920 1.120 ;
 END
END CK
PIN A0
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 107.320 0.000 108.440 1.120 ;
  LAYER ME3 ;
  RECT 107.320 0.000 108.440 1.120 ;
  LAYER ME2 ;
  RECT 107.320 0.000 108.440 1.120 ;
  LAYER ME1 ;
  RECT 107.320 0.000 108.440 1.120 ;
 END
END A0
PIN A3
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 102.980 0.000 104.100 1.120 ;
  LAYER ME3 ;
  RECT 102.980 0.000 104.100 1.120 ;
  LAYER ME2 ;
  RECT 102.980 0.000 104.100 1.120 ;
  LAYER ME1 ;
  RECT 102.980 0.000 104.100 1.120 ;
 END
END A3
PIN A4
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 95.540 0.000 96.660 1.120 ;
  LAYER ME3 ;
  RECT 95.540 0.000 96.660 1.120 ;
  LAYER ME2 ;
  RECT 95.540 0.000 96.660 1.120 ;
  LAYER ME1 ;
  RECT 95.540 0.000 96.660 1.120 ;
 END
END A4
PIN A5
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 92.440 0.000 93.560 1.120 ;
  LAYER ME3 ;
  RECT 92.440 0.000 93.560 1.120 ;
  LAYER ME2 ;
  RECT 92.440 0.000 93.560 1.120 ;
  LAYER ME1 ;
  RECT 92.440 0.000 93.560 1.120 ;
 END
END A5
PIN A6
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 85.000 0.000 86.120 1.120 ;
  LAYER ME3 ;
  RECT 85.000 0.000 86.120 1.120 ;
  LAYER ME2 ;
  RECT 85.000 0.000 86.120 1.120 ;
  LAYER ME1 ;
  RECT 85.000 0.000 86.120 1.120 ;
 END
END A6
PIN A7
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 81.900 0.000 83.020 1.120 ;
  LAYER ME3 ;
  RECT 81.900 0.000 83.020 1.120 ;
  LAYER ME2 ;
  RECT 81.900 0.000 83.020 1.120 ;
  LAYER ME1 ;
  RECT 81.900 0.000 83.020 1.120 ;
 END
END A7
PIN A8
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 74.460 0.000 75.580 1.120 ;
  LAYER ME3 ;
  RECT 74.460 0.000 75.580 1.120 ;
  LAYER ME2 ;
  RECT 74.460 0.000 75.580 1.120 ;
  LAYER ME1 ;
  RECT 74.460 0.000 75.580 1.120 ;
 END
END A8
PIN DO3
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 63.300 0.000 64.420 1.120 ;
  LAYER ME3 ;
  RECT 63.300 0.000 64.420 1.120 ;
  LAYER ME2 ;
  RECT 63.300 0.000 64.420 1.120 ;
  LAYER ME1 ;
  RECT 63.300 0.000 64.420 1.120 ;
 END
END DO3
PIN DI3
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 54.620 0.000 55.740 1.120 ;
  LAYER ME3 ;
  RECT 54.620 0.000 55.740 1.120 ;
  LAYER ME2 ;
  RECT 54.620 0.000 55.740 1.120 ;
  LAYER ME1 ;
  RECT 54.620 0.000 55.740 1.120 ;
 END
END DI3
PIN DO2
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 50.280 0.000 51.400 1.120 ;
  LAYER ME3 ;
  RECT 50.280 0.000 51.400 1.120 ;
  LAYER ME2 ;
  RECT 50.280 0.000 51.400 1.120 ;
  LAYER ME1 ;
  RECT 50.280 0.000 51.400 1.120 ;
 END
END DO2
PIN DI2
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 41.600 0.000 42.720 1.120 ;
  LAYER ME3 ;
  RECT 41.600 0.000 42.720 1.120 ;
  LAYER ME2 ;
  RECT 41.600 0.000 42.720 1.120 ;
  LAYER ME1 ;
  RECT 41.600 0.000 42.720 1.120 ;
 END
END DI2
PIN DO1
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 33.540 0.000 34.660 1.120 ;
  LAYER ME3 ;
  RECT 33.540 0.000 34.660 1.120 ;
  LAYER ME2 ;
  RECT 33.540 0.000 34.660 1.120 ;
  LAYER ME1 ;
  RECT 33.540 0.000 34.660 1.120 ;
 END
END DO1
PIN DI1
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 24.860 0.000 25.980 1.120 ;
  LAYER ME3 ;
  RECT 24.860 0.000 25.980 1.120 ;
  LAYER ME2 ;
  RECT 24.860 0.000 25.980 1.120 ;
  LAYER ME1 ;
  RECT 24.860 0.000 25.980 1.120 ;
 END
END DI1
PIN DO0
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 19.900 0.000 21.020 1.120 ;
  LAYER ME3 ;
  RECT 19.900 0.000 21.020 1.120 ;
  LAYER ME2 ;
  RECT 19.900 0.000 21.020 1.120 ;
  LAYER ME1 ;
  RECT 19.900 0.000 21.020 1.120 ;
 END
END DO0
PIN DI0
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 11.840 0.000 12.960 1.120 ;
  LAYER ME3 ;
  RECT 11.840 0.000 12.960 1.120 ;
  LAYER ME2 ;
  RECT 11.840 0.000 12.960 1.120 ;
  LAYER ME1 ;
  RECT 11.840 0.000 12.960 1.120 ;
 END
END DI0
OBS
  LAYER ME1 SPACING 0.280 ;
  RECT 0.000 0.140 213.900 259.840 ;
  LAYER ME2 SPACING 0.320 ;
  RECT 0.000 0.140 213.900 259.840 ;
  LAYER ME3 SPACING 0.320 ;
  RECT 0.000 0.140 213.900 259.840 ;
  LAYER ME4 SPACING 0.600 ;
  RECT 0.000 0.140 213.900 259.840 ;
  LAYER VI1 ;
  RECT 0.000 0.140 213.900 259.840 ;
  LAYER VI2 ;
  RECT 0.000 0.140 213.900 259.840 ;
  LAYER VI3 ;
  RECT 0.000 0.140 213.900 259.840 ;
END
END SUMA_400_M1
END LIBRARY



