# 
#              Synchronous High Speed Single Port SRAM Compiler 
# 
#                    UMC 0.18um GenericII Logic Process
#    __________________________________________________________________________
# 
# 
#      (C) Copyright 2002-2009 Faraday Technology Corp. All Rights Reserved.
#    
#    This source code is an unpublished work belongs to Faraday Technology
#    Corp.  It is considered a trade secret and is not to be divulged or
#    used by parties who have not received written authorization from
#    Faraday Technology Corp.
#    
#    Faraday's home page can be found at:
#    http://www.faraday-tech.com/
#   
#       Module Name      : SUMA_1296
#       Words            : 1296
#       Bits             : 20
#       Byte-Write       : 1
#       Aspect Ratio     : 1
#       Output Loading   : 0.05  (pf)
#       Data Slew        : 0.02  (ns)
#       CK Slew          : 0.02  (ns)
#       Power Ring Width : 2  (um)
# 
# -----------------------------------------------------------------------------
# 
#       Library          : FSA0M_A
#       Memaker          : 200901.2.1
#       Date             : 2024/03/30 23:44:28
# 
# -----------------------------------------------------------------------------


NAMESCASESENSITIVE ON ;
MACRO SUMA_1296
CLASS BLOCK ;
FOREIGN SUMA_1296 0.000 0.000 ;
ORIGIN 0.000 0.000 ;
SIZE 397.420 BY 534.240 ;
SYMMETRY x y r90 ;
SITE core ;
PIN GND
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
 PORT
  LAYER ME4 ;
  RECT 396.300 521.700 397.420 524.940 ;
  LAYER ME3 ;
  RECT 396.300 521.700 397.420 524.940 ;
  LAYER ME2 ;
  RECT 396.300 521.700 397.420 524.940 ;
  LAYER ME1 ;
  RECT 396.300 521.700 397.420 524.940 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 513.860 397.420 517.100 ;
  LAYER ME3 ;
  RECT 396.300 513.860 397.420 517.100 ;
  LAYER ME2 ;
  RECT 396.300 513.860 397.420 517.100 ;
  LAYER ME1 ;
  RECT 396.300 513.860 397.420 517.100 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 506.020 397.420 509.260 ;
  LAYER ME3 ;
  RECT 396.300 506.020 397.420 509.260 ;
  LAYER ME2 ;
  RECT 396.300 506.020 397.420 509.260 ;
  LAYER ME1 ;
  RECT 396.300 506.020 397.420 509.260 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 498.180 397.420 501.420 ;
  LAYER ME3 ;
  RECT 396.300 498.180 397.420 501.420 ;
  LAYER ME2 ;
  RECT 396.300 498.180 397.420 501.420 ;
  LAYER ME1 ;
  RECT 396.300 498.180 397.420 501.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 490.340 397.420 493.580 ;
  LAYER ME3 ;
  RECT 396.300 490.340 397.420 493.580 ;
  LAYER ME2 ;
  RECT 396.300 490.340 397.420 493.580 ;
  LAYER ME1 ;
  RECT 396.300 490.340 397.420 493.580 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 482.500 397.420 485.740 ;
  LAYER ME3 ;
  RECT 396.300 482.500 397.420 485.740 ;
  LAYER ME2 ;
  RECT 396.300 482.500 397.420 485.740 ;
  LAYER ME1 ;
  RECT 396.300 482.500 397.420 485.740 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 443.300 397.420 446.540 ;
  LAYER ME3 ;
  RECT 396.300 443.300 397.420 446.540 ;
  LAYER ME2 ;
  RECT 396.300 443.300 397.420 446.540 ;
  LAYER ME1 ;
  RECT 396.300 443.300 397.420 446.540 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 435.460 397.420 438.700 ;
  LAYER ME3 ;
  RECT 396.300 435.460 397.420 438.700 ;
  LAYER ME2 ;
  RECT 396.300 435.460 397.420 438.700 ;
  LAYER ME1 ;
  RECT 396.300 435.460 397.420 438.700 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 427.620 397.420 430.860 ;
  LAYER ME3 ;
  RECT 396.300 427.620 397.420 430.860 ;
  LAYER ME2 ;
  RECT 396.300 427.620 397.420 430.860 ;
  LAYER ME1 ;
  RECT 396.300 427.620 397.420 430.860 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 419.780 397.420 423.020 ;
  LAYER ME3 ;
  RECT 396.300 419.780 397.420 423.020 ;
  LAYER ME2 ;
  RECT 396.300 419.780 397.420 423.020 ;
  LAYER ME1 ;
  RECT 396.300 419.780 397.420 423.020 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 411.940 397.420 415.180 ;
  LAYER ME3 ;
  RECT 396.300 411.940 397.420 415.180 ;
  LAYER ME2 ;
  RECT 396.300 411.940 397.420 415.180 ;
  LAYER ME1 ;
  RECT 396.300 411.940 397.420 415.180 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 404.100 397.420 407.340 ;
  LAYER ME3 ;
  RECT 396.300 404.100 397.420 407.340 ;
  LAYER ME2 ;
  RECT 396.300 404.100 397.420 407.340 ;
  LAYER ME1 ;
  RECT 396.300 404.100 397.420 407.340 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 364.900 397.420 368.140 ;
  LAYER ME3 ;
  RECT 396.300 364.900 397.420 368.140 ;
  LAYER ME2 ;
  RECT 396.300 364.900 397.420 368.140 ;
  LAYER ME1 ;
  RECT 396.300 364.900 397.420 368.140 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 357.060 397.420 360.300 ;
  LAYER ME3 ;
  RECT 396.300 357.060 397.420 360.300 ;
  LAYER ME2 ;
  RECT 396.300 357.060 397.420 360.300 ;
  LAYER ME1 ;
  RECT 396.300 357.060 397.420 360.300 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 349.220 397.420 352.460 ;
  LAYER ME3 ;
  RECT 396.300 349.220 397.420 352.460 ;
  LAYER ME2 ;
  RECT 396.300 349.220 397.420 352.460 ;
  LAYER ME1 ;
  RECT 396.300 349.220 397.420 352.460 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 341.380 397.420 344.620 ;
  LAYER ME3 ;
  RECT 396.300 341.380 397.420 344.620 ;
  LAYER ME2 ;
  RECT 396.300 341.380 397.420 344.620 ;
  LAYER ME1 ;
  RECT 396.300 341.380 397.420 344.620 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 333.540 397.420 336.780 ;
  LAYER ME3 ;
  RECT 396.300 333.540 397.420 336.780 ;
  LAYER ME2 ;
  RECT 396.300 333.540 397.420 336.780 ;
  LAYER ME1 ;
  RECT 396.300 333.540 397.420 336.780 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 325.700 397.420 328.940 ;
  LAYER ME3 ;
  RECT 396.300 325.700 397.420 328.940 ;
  LAYER ME2 ;
  RECT 396.300 325.700 397.420 328.940 ;
  LAYER ME1 ;
  RECT 396.300 325.700 397.420 328.940 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 286.500 397.420 289.740 ;
  LAYER ME3 ;
  RECT 396.300 286.500 397.420 289.740 ;
  LAYER ME2 ;
  RECT 396.300 286.500 397.420 289.740 ;
  LAYER ME1 ;
  RECT 396.300 286.500 397.420 289.740 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 278.660 397.420 281.900 ;
  LAYER ME3 ;
  RECT 396.300 278.660 397.420 281.900 ;
  LAYER ME2 ;
  RECT 396.300 278.660 397.420 281.900 ;
  LAYER ME1 ;
  RECT 396.300 278.660 397.420 281.900 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 270.820 397.420 274.060 ;
  LAYER ME3 ;
  RECT 396.300 270.820 397.420 274.060 ;
  LAYER ME2 ;
  RECT 396.300 270.820 397.420 274.060 ;
  LAYER ME1 ;
  RECT 396.300 270.820 397.420 274.060 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 262.980 397.420 266.220 ;
  LAYER ME3 ;
  RECT 396.300 262.980 397.420 266.220 ;
  LAYER ME2 ;
  RECT 396.300 262.980 397.420 266.220 ;
  LAYER ME1 ;
  RECT 396.300 262.980 397.420 266.220 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 255.140 397.420 258.380 ;
  LAYER ME3 ;
  RECT 396.300 255.140 397.420 258.380 ;
  LAYER ME2 ;
  RECT 396.300 255.140 397.420 258.380 ;
  LAYER ME1 ;
  RECT 396.300 255.140 397.420 258.380 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 247.300 397.420 250.540 ;
  LAYER ME3 ;
  RECT 396.300 247.300 397.420 250.540 ;
  LAYER ME2 ;
  RECT 396.300 247.300 397.420 250.540 ;
  LAYER ME1 ;
  RECT 396.300 247.300 397.420 250.540 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 208.100 397.420 211.340 ;
  LAYER ME3 ;
  RECT 396.300 208.100 397.420 211.340 ;
  LAYER ME2 ;
  RECT 396.300 208.100 397.420 211.340 ;
  LAYER ME1 ;
  RECT 396.300 208.100 397.420 211.340 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 200.260 397.420 203.500 ;
  LAYER ME3 ;
  RECT 396.300 200.260 397.420 203.500 ;
  LAYER ME2 ;
  RECT 396.300 200.260 397.420 203.500 ;
  LAYER ME1 ;
  RECT 396.300 200.260 397.420 203.500 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 192.420 397.420 195.660 ;
  LAYER ME3 ;
  RECT 396.300 192.420 397.420 195.660 ;
  LAYER ME2 ;
  RECT 396.300 192.420 397.420 195.660 ;
  LAYER ME1 ;
  RECT 396.300 192.420 397.420 195.660 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 184.580 397.420 187.820 ;
  LAYER ME3 ;
  RECT 396.300 184.580 397.420 187.820 ;
  LAYER ME2 ;
  RECT 396.300 184.580 397.420 187.820 ;
  LAYER ME1 ;
  RECT 396.300 184.580 397.420 187.820 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 176.740 397.420 179.980 ;
  LAYER ME3 ;
  RECT 396.300 176.740 397.420 179.980 ;
  LAYER ME2 ;
  RECT 396.300 176.740 397.420 179.980 ;
  LAYER ME1 ;
  RECT 396.300 176.740 397.420 179.980 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 168.900 397.420 172.140 ;
  LAYER ME3 ;
  RECT 396.300 168.900 397.420 172.140 ;
  LAYER ME2 ;
  RECT 396.300 168.900 397.420 172.140 ;
  LAYER ME1 ;
  RECT 396.300 168.900 397.420 172.140 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 129.700 397.420 132.940 ;
  LAYER ME3 ;
  RECT 396.300 129.700 397.420 132.940 ;
  LAYER ME2 ;
  RECT 396.300 129.700 397.420 132.940 ;
  LAYER ME1 ;
  RECT 396.300 129.700 397.420 132.940 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 121.860 397.420 125.100 ;
  LAYER ME3 ;
  RECT 396.300 121.860 397.420 125.100 ;
  LAYER ME2 ;
  RECT 396.300 121.860 397.420 125.100 ;
  LAYER ME1 ;
  RECT 396.300 121.860 397.420 125.100 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 114.020 397.420 117.260 ;
  LAYER ME3 ;
  RECT 396.300 114.020 397.420 117.260 ;
  LAYER ME2 ;
  RECT 396.300 114.020 397.420 117.260 ;
  LAYER ME1 ;
  RECT 396.300 114.020 397.420 117.260 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 106.180 397.420 109.420 ;
  LAYER ME3 ;
  RECT 396.300 106.180 397.420 109.420 ;
  LAYER ME2 ;
  RECT 396.300 106.180 397.420 109.420 ;
  LAYER ME1 ;
  RECT 396.300 106.180 397.420 109.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 98.340 397.420 101.580 ;
  LAYER ME3 ;
  RECT 396.300 98.340 397.420 101.580 ;
  LAYER ME2 ;
  RECT 396.300 98.340 397.420 101.580 ;
  LAYER ME1 ;
  RECT 396.300 98.340 397.420 101.580 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 90.500 397.420 93.740 ;
  LAYER ME3 ;
  RECT 396.300 90.500 397.420 93.740 ;
  LAYER ME2 ;
  RECT 396.300 90.500 397.420 93.740 ;
  LAYER ME1 ;
  RECT 396.300 90.500 397.420 93.740 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 51.300 397.420 54.540 ;
  LAYER ME3 ;
  RECT 396.300 51.300 397.420 54.540 ;
  LAYER ME2 ;
  RECT 396.300 51.300 397.420 54.540 ;
  LAYER ME1 ;
  RECT 396.300 51.300 397.420 54.540 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 43.460 397.420 46.700 ;
  LAYER ME3 ;
  RECT 396.300 43.460 397.420 46.700 ;
  LAYER ME2 ;
  RECT 396.300 43.460 397.420 46.700 ;
  LAYER ME1 ;
  RECT 396.300 43.460 397.420 46.700 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 35.620 397.420 38.860 ;
  LAYER ME3 ;
  RECT 396.300 35.620 397.420 38.860 ;
  LAYER ME2 ;
  RECT 396.300 35.620 397.420 38.860 ;
  LAYER ME1 ;
  RECT 396.300 35.620 397.420 38.860 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 27.780 397.420 31.020 ;
  LAYER ME3 ;
  RECT 396.300 27.780 397.420 31.020 ;
  LAYER ME2 ;
  RECT 396.300 27.780 397.420 31.020 ;
  LAYER ME1 ;
  RECT 396.300 27.780 397.420 31.020 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 19.940 397.420 23.180 ;
  LAYER ME3 ;
  RECT 396.300 19.940 397.420 23.180 ;
  LAYER ME2 ;
  RECT 396.300 19.940 397.420 23.180 ;
  LAYER ME1 ;
  RECT 396.300 19.940 397.420 23.180 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 12.100 397.420 15.340 ;
  LAYER ME3 ;
  RECT 396.300 12.100 397.420 15.340 ;
  LAYER ME2 ;
  RECT 396.300 12.100 397.420 15.340 ;
  LAYER ME1 ;
  RECT 396.300 12.100 397.420 15.340 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 521.700 1.120 524.940 ;
  LAYER ME3 ;
  RECT 0.000 521.700 1.120 524.940 ;
  LAYER ME2 ;
  RECT 0.000 521.700 1.120 524.940 ;
  LAYER ME1 ;
  RECT 0.000 521.700 1.120 524.940 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 513.860 1.120 517.100 ;
  LAYER ME3 ;
  RECT 0.000 513.860 1.120 517.100 ;
  LAYER ME2 ;
  RECT 0.000 513.860 1.120 517.100 ;
  LAYER ME1 ;
  RECT 0.000 513.860 1.120 517.100 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 506.020 1.120 509.260 ;
  LAYER ME3 ;
  RECT 0.000 506.020 1.120 509.260 ;
  LAYER ME2 ;
  RECT 0.000 506.020 1.120 509.260 ;
  LAYER ME1 ;
  RECT 0.000 506.020 1.120 509.260 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 498.180 1.120 501.420 ;
  LAYER ME3 ;
  RECT 0.000 498.180 1.120 501.420 ;
  LAYER ME2 ;
  RECT 0.000 498.180 1.120 501.420 ;
  LAYER ME1 ;
  RECT 0.000 498.180 1.120 501.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 490.340 1.120 493.580 ;
  LAYER ME3 ;
  RECT 0.000 490.340 1.120 493.580 ;
  LAYER ME2 ;
  RECT 0.000 490.340 1.120 493.580 ;
  LAYER ME1 ;
  RECT 0.000 490.340 1.120 493.580 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 482.500 1.120 485.740 ;
  LAYER ME3 ;
  RECT 0.000 482.500 1.120 485.740 ;
  LAYER ME2 ;
  RECT 0.000 482.500 1.120 485.740 ;
  LAYER ME1 ;
  RECT 0.000 482.500 1.120 485.740 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 443.300 1.120 446.540 ;
  LAYER ME3 ;
  RECT 0.000 443.300 1.120 446.540 ;
  LAYER ME2 ;
  RECT 0.000 443.300 1.120 446.540 ;
  LAYER ME1 ;
  RECT 0.000 443.300 1.120 446.540 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 435.460 1.120 438.700 ;
  LAYER ME3 ;
  RECT 0.000 435.460 1.120 438.700 ;
  LAYER ME2 ;
  RECT 0.000 435.460 1.120 438.700 ;
  LAYER ME1 ;
  RECT 0.000 435.460 1.120 438.700 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 427.620 1.120 430.860 ;
  LAYER ME3 ;
  RECT 0.000 427.620 1.120 430.860 ;
  LAYER ME2 ;
  RECT 0.000 427.620 1.120 430.860 ;
  LAYER ME1 ;
  RECT 0.000 427.620 1.120 430.860 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 419.780 1.120 423.020 ;
  LAYER ME3 ;
  RECT 0.000 419.780 1.120 423.020 ;
  LAYER ME2 ;
  RECT 0.000 419.780 1.120 423.020 ;
  LAYER ME1 ;
  RECT 0.000 419.780 1.120 423.020 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 411.940 1.120 415.180 ;
  LAYER ME3 ;
  RECT 0.000 411.940 1.120 415.180 ;
  LAYER ME2 ;
  RECT 0.000 411.940 1.120 415.180 ;
  LAYER ME1 ;
  RECT 0.000 411.940 1.120 415.180 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 404.100 1.120 407.340 ;
  LAYER ME3 ;
  RECT 0.000 404.100 1.120 407.340 ;
  LAYER ME2 ;
  RECT 0.000 404.100 1.120 407.340 ;
  LAYER ME1 ;
  RECT 0.000 404.100 1.120 407.340 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 364.900 1.120 368.140 ;
  LAYER ME3 ;
  RECT 0.000 364.900 1.120 368.140 ;
  LAYER ME2 ;
  RECT 0.000 364.900 1.120 368.140 ;
  LAYER ME1 ;
  RECT 0.000 364.900 1.120 368.140 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 357.060 1.120 360.300 ;
  LAYER ME3 ;
  RECT 0.000 357.060 1.120 360.300 ;
  LAYER ME2 ;
  RECT 0.000 357.060 1.120 360.300 ;
  LAYER ME1 ;
  RECT 0.000 357.060 1.120 360.300 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 349.220 1.120 352.460 ;
  LAYER ME3 ;
  RECT 0.000 349.220 1.120 352.460 ;
  LAYER ME2 ;
  RECT 0.000 349.220 1.120 352.460 ;
  LAYER ME1 ;
  RECT 0.000 349.220 1.120 352.460 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 341.380 1.120 344.620 ;
  LAYER ME3 ;
  RECT 0.000 341.380 1.120 344.620 ;
  LAYER ME2 ;
  RECT 0.000 341.380 1.120 344.620 ;
  LAYER ME1 ;
  RECT 0.000 341.380 1.120 344.620 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 333.540 1.120 336.780 ;
  LAYER ME3 ;
  RECT 0.000 333.540 1.120 336.780 ;
  LAYER ME2 ;
  RECT 0.000 333.540 1.120 336.780 ;
  LAYER ME1 ;
  RECT 0.000 333.540 1.120 336.780 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 325.700 1.120 328.940 ;
  LAYER ME3 ;
  RECT 0.000 325.700 1.120 328.940 ;
  LAYER ME2 ;
  RECT 0.000 325.700 1.120 328.940 ;
  LAYER ME1 ;
  RECT 0.000 325.700 1.120 328.940 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 286.500 1.120 289.740 ;
  LAYER ME3 ;
  RECT 0.000 286.500 1.120 289.740 ;
  LAYER ME2 ;
  RECT 0.000 286.500 1.120 289.740 ;
  LAYER ME1 ;
  RECT 0.000 286.500 1.120 289.740 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 278.660 1.120 281.900 ;
  LAYER ME3 ;
  RECT 0.000 278.660 1.120 281.900 ;
  LAYER ME2 ;
  RECT 0.000 278.660 1.120 281.900 ;
  LAYER ME1 ;
  RECT 0.000 278.660 1.120 281.900 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 270.820 1.120 274.060 ;
  LAYER ME3 ;
  RECT 0.000 270.820 1.120 274.060 ;
  LAYER ME2 ;
  RECT 0.000 270.820 1.120 274.060 ;
  LAYER ME1 ;
  RECT 0.000 270.820 1.120 274.060 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 262.980 1.120 266.220 ;
  LAYER ME3 ;
  RECT 0.000 262.980 1.120 266.220 ;
  LAYER ME2 ;
  RECT 0.000 262.980 1.120 266.220 ;
  LAYER ME1 ;
  RECT 0.000 262.980 1.120 266.220 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 255.140 1.120 258.380 ;
  LAYER ME3 ;
  RECT 0.000 255.140 1.120 258.380 ;
  LAYER ME2 ;
  RECT 0.000 255.140 1.120 258.380 ;
  LAYER ME1 ;
  RECT 0.000 255.140 1.120 258.380 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 247.300 1.120 250.540 ;
  LAYER ME3 ;
  RECT 0.000 247.300 1.120 250.540 ;
  LAYER ME2 ;
  RECT 0.000 247.300 1.120 250.540 ;
  LAYER ME1 ;
  RECT 0.000 247.300 1.120 250.540 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 208.100 1.120 211.340 ;
  LAYER ME3 ;
  RECT 0.000 208.100 1.120 211.340 ;
  LAYER ME2 ;
  RECT 0.000 208.100 1.120 211.340 ;
  LAYER ME1 ;
  RECT 0.000 208.100 1.120 211.340 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 200.260 1.120 203.500 ;
  LAYER ME3 ;
  RECT 0.000 200.260 1.120 203.500 ;
  LAYER ME2 ;
  RECT 0.000 200.260 1.120 203.500 ;
  LAYER ME1 ;
  RECT 0.000 200.260 1.120 203.500 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 192.420 1.120 195.660 ;
  LAYER ME3 ;
  RECT 0.000 192.420 1.120 195.660 ;
  LAYER ME2 ;
  RECT 0.000 192.420 1.120 195.660 ;
  LAYER ME1 ;
  RECT 0.000 192.420 1.120 195.660 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 184.580 1.120 187.820 ;
  LAYER ME3 ;
  RECT 0.000 184.580 1.120 187.820 ;
  LAYER ME2 ;
  RECT 0.000 184.580 1.120 187.820 ;
  LAYER ME1 ;
  RECT 0.000 184.580 1.120 187.820 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 176.740 1.120 179.980 ;
  LAYER ME3 ;
  RECT 0.000 176.740 1.120 179.980 ;
  LAYER ME2 ;
  RECT 0.000 176.740 1.120 179.980 ;
  LAYER ME1 ;
  RECT 0.000 176.740 1.120 179.980 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 168.900 1.120 172.140 ;
  LAYER ME3 ;
  RECT 0.000 168.900 1.120 172.140 ;
  LAYER ME2 ;
  RECT 0.000 168.900 1.120 172.140 ;
  LAYER ME1 ;
  RECT 0.000 168.900 1.120 172.140 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 129.700 1.120 132.940 ;
  LAYER ME3 ;
  RECT 0.000 129.700 1.120 132.940 ;
  LAYER ME2 ;
  RECT 0.000 129.700 1.120 132.940 ;
  LAYER ME1 ;
  RECT 0.000 129.700 1.120 132.940 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 121.860 1.120 125.100 ;
  LAYER ME3 ;
  RECT 0.000 121.860 1.120 125.100 ;
  LAYER ME2 ;
  RECT 0.000 121.860 1.120 125.100 ;
  LAYER ME1 ;
  RECT 0.000 121.860 1.120 125.100 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 114.020 1.120 117.260 ;
  LAYER ME3 ;
  RECT 0.000 114.020 1.120 117.260 ;
  LAYER ME2 ;
  RECT 0.000 114.020 1.120 117.260 ;
  LAYER ME1 ;
  RECT 0.000 114.020 1.120 117.260 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 106.180 1.120 109.420 ;
  LAYER ME3 ;
  RECT 0.000 106.180 1.120 109.420 ;
  LAYER ME2 ;
  RECT 0.000 106.180 1.120 109.420 ;
  LAYER ME1 ;
  RECT 0.000 106.180 1.120 109.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 98.340 1.120 101.580 ;
  LAYER ME3 ;
  RECT 0.000 98.340 1.120 101.580 ;
  LAYER ME2 ;
  RECT 0.000 98.340 1.120 101.580 ;
  LAYER ME1 ;
  RECT 0.000 98.340 1.120 101.580 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 90.500 1.120 93.740 ;
  LAYER ME3 ;
  RECT 0.000 90.500 1.120 93.740 ;
  LAYER ME2 ;
  RECT 0.000 90.500 1.120 93.740 ;
  LAYER ME1 ;
  RECT 0.000 90.500 1.120 93.740 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 51.300 1.120 54.540 ;
  LAYER ME3 ;
  RECT 0.000 51.300 1.120 54.540 ;
  LAYER ME2 ;
  RECT 0.000 51.300 1.120 54.540 ;
  LAYER ME1 ;
  RECT 0.000 51.300 1.120 54.540 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 43.460 1.120 46.700 ;
  LAYER ME3 ;
  RECT 0.000 43.460 1.120 46.700 ;
  LAYER ME2 ;
  RECT 0.000 43.460 1.120 46.700 ;
  LAYER ME1 ;
  RECT 0.000 43.460 1.120 46.700 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 35.620 1.120 38.860 ;
  LAYER ME3 ;
  RECT 0.000 35.620 1.120 38.860 ;
  LAYER ME2 ;
  RECT 0.000 35.620 1.120 38.860 ;
  LAYER ME1 ;
  RECT 0.000 35.620 1.120 38.860 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 27.780 1.120 31.020 ;
  LAYER ME3 ;
  RECT 0.000 27.780 1.120 31.020 ;
  LAYER ME2 ;
  RECT 0.000 27.780 1.120 31.020 ;
  LAYER ME1 ;
  RECT 0.000 27.780 1.120 31.020 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 19.940 1.120 23.180 ;
  LAYER ME3 ;
  RECT 0.000 19.940 1.120 23.180 ;
  LAYER ME2 ;
  RECT 0.000 19.940 1.120 23.180 ;
  LAYER ME1 ;
  RECT 0.000 19.940 1.120 23.180 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 12.100 1.120 15.340 ;
  LAYER ME3 ;
  RECT 0.000 12.100 1.120 15.340 ;
  LAYER ME2 ;
  RECT 0.000 12.100 1.120 15.340 ;
  LAYER ME1 ;
  RECT 0.000 12.100 1.120 15.340 ;
 END
 PORT
  LAYER ME4 ;
  RECT 385.420 533.120 388.960 534.240 ;
  LAYER ME3 ;
  RECT 385.420 533.120 388.960 534.240 ;
  LAYER ME2 ;
  RECT 385.420 533.120 388.960 534.240 ;
  LAYER ME1 ;
  RECT 385.420 533.120 388.960 534.240 ;
 END
 PORT
  LAYER ME4 ;
  RECT 376.740 533.120 380.280 534.240 ;
  LAYER ME3 ;
  RECT 376.740 533.120 380.280 534.240 ;
  LAYER ME2 ;
  RECT 376.740 533.120 380.280 534.240 ;
  LAYER ME1 ;
  RECT 376.740 533.120 380.280 534.240 ;
 END
 PORT
  LAYER ME4 ;
  RECT 368.060 533.120 371.600 534.240 ;
  LAYER ME3 ;
  RECT 368.060 533.120 371.600 534.240 ;
  LAYER ME2 ;
  RECT 368.060 533.120 371.600 534.240 ;
  LAYER ME1 ;
  RECT 368.060 533.120 371.600 534.240 ;
 END
 PORT
  LAYER ME4 ;
  RECT 359.380 533.120 362.920 534.240 ;
  LAYER ME3 ;
  RECT 359.380 533.120 362.920 534.240 ;
  LAYER ME2 ;
  RECT 359.380 533.120 362.920 534.240 ;
  LAYER ME1 ;
  RECT 359.380 533.120 362.920 534.240 ;
 END
 PORT
  LAYER ME4 ;
  RECT 315.980 533.120 319.520 534.240 ;
  LAYER ME3 ;
  RECT 315.980 533.120 319.520 534.240 ;
  LAYER ME2 ;
  RECT 315.980 533.120 319.520 534.240 ;
  LAYER ME1 ;
  RECT 315.980 533.120 319.520 534.240 ;
 END
 PORT
  LAYER ME4 ;
  RECT 307.300 533.120 310.840 534.240 ;
  LAYER ME3 ;
  RECT 307.300 533.120 310.840 534.240 ;
  LAYER ME2 ;
  RECT 307.300 533.120 310.840 534.240 ;
  LAYER ME1 ;
  RECT 307.300 533.120 310.840 534.240 ;
 END
 PORT
  LAYER ME4 ;
  RECT 298.620 533.120 302.160 534.240 ;
  LAYER ME3 ;
  RECT 298.620 533.120 302.160 534.240 ;
  LAYER ME2 ;
  RECT 298.620 533.120 302.160 534.240 ;
  LAYER ME1 ;
  RECT 298.620 533.120 302.160 534.240 ;
 END
 PORT
  LAYER ME4 ;
  RECT 289.940 533.120 293.480 534.240 ;
  LAYER ME3 ;
  RECT 289.940 533.120 293.480 534.240 ;
  LAYER ME2 ;
  RECT 289.940 533.120 293.480 534.240 ;
  LAYER ME1 ;
  RECT 289.940 533.120 293.480 534.240 ;
 END
 PORT
  LAYER ME4 ;
  RECT 281.260 533.120 284.800 534.240 ;
  LAYER ME3 ;
  RECT 281.260 533.120 284.800 534.240 ;
  LAYER ME2 ;
  RECT 281.260 533.120 284.800 534.240 ;
  LAYER ME1 ;
  RECT 281.260 533.120 284.800 534.240 ;
 END
 PORT
  LAYER ME4 ;
  RECT 272.580 533.120 276.120 534.240 ;
  LAYER ME3 ;
  RECT 272.580 533.120 276.120 534.240 ;
  LAYER ME2 ;
  RECT 272.580 533.120 276.120 534.240 ;
  LAYER ME1 ;
  RECT 272.580 533.120 276.120 534.240 ;
 END
 PORT
  LAYER ME4 ;
  RECT 229.180 533.120 232.720 534.240 ;
  LAYER ME3 ;
  RECT 229.180 533.120 232.720 534.240 ;
  LAYER ME2 ;
  RECT 229.180 533.120 232.720 534.240 ;
  LAYER ME1 ;
  RECT 229.180 533.120 232.720 534.240 ;
 END
 PORT
  LAYER ME4 ;
  RECT 220.500 533.120 224.040 534.240 ;
  LAYER ME3 ;
  RECT 220.500 533.120 224.040 534.240 ;
  LAYER ME2 ;
  RECT 220.500 533.120 224.040 534.240 ;
  LAYER ME1 ;
  RECT 220.500 533.120 224.040 534.240 ;
 END
 PORT
  LAYER ME4 ;
  RECT 211.820 533.120 215.360 534.240 ;
  LAYER ME3 ;
  RECT 211.820 533.120 215.360 534.240 ;
  LAYER ME2 ;
  RECT 211.820 533.120 215.360 534.240 ;
  LAYER ME1 ;
  RECT 211.820 533.120 215.360 534.240 ;
 END
 PORT
  LAYER ME4 ;
  RECT 203.140 533.120 206.680 534.240 ;
  LAYER ME3 ;
  RECT 203.140 533.120 206.680 534.240 ;
  LAYER ME2 ;
  RECT 203.140 533.120 206.680 534.240 ;
  LAYER ME1 ;
  RECT 203.140 533.120 206.680 534.240 ;
 END
 PORT
  LAYER ME4 ;
  RECT 194.460 533.120 198.000 534.240 ;
  LAYER ME3 ;
  RECT 194.460 533.120 198.000 534.240 ;
  LAYER ME2 ;
  RECT 194.460 533.120 198.000 534.240 ;
  LAYER ME1 ;
  RECT 194.460 533.120 198.000 534.240 ;
 END
 PORT
  LAYER ME4 ;
  RECT 185.780 533.120 189.320 534.240 ;
  LAYER ME3 ;
  RECT 185.780 533.120 189.320 534.240 ;
  LAYER ME2 ;
  RECT 185.780 533.120 189.320 534.240 ;
  LAYER ME1 ;
  RECT 185.780 533.120 189.320 534.240 ;
 END
 PORT
  LAYER ME4 ;
  RECT 142.380 533.120 145.920 534.240 ;
  LAYER ME3 ;
  RECT 142.380 533.120 145.920 534.240 ;
  LAYER ME2 ;
  RECT 142.380 533.120 145.920 534.240 ;
  LAYER ME1 ;
  RECT 142.380 533.120 145.920 534.240 ;
 END
 PORT
  LAYER ME4 ;
  RECT 133.700 533.120 137.240 534.240 ;
  LAYER ME3 ;
  RECT 133.700 533.120 137.240 534.240 ;
  LAYER ME2 ;
  RECT 133.700 533.120 137.240 534.240 ;
  LAYER ME1 ;
  RECT 133.700 533.120 137.240 534.240 ;
 END
 PORT
  LAYER ME4 ;
  RECT 125.020 533.120 128.560 534.240 ;
  LAYER ME3 ;
  RECT 125.020 533.120 128.560 534.240 ;
  LAYER ME2 ;
  RECT 125.020 533.120 128.560 534.240 ;
  LAYER ME1 ;
  RECT 125.020 533.120 128.560 534.240 ;
 END
 PORT
  LAYER ME4 ;
  RECT 116.340 533.120 119.880 534.240 ;
  LAYER ME3 ;
  RECT 116.340 533.120 119.880 534.240 ;
  LAYER ME2 ;
  RECT 116.340 533.120 119.880 534.240 ;
  LAYER ME1 ;
  RECT 116.340 533.120 119.880 534.240 ;
 END
 PORT
  LAYER ME4 ;
  RECT 107.660 533.120 111.200 534.240 ;
  LAYER ME3 ;
  RECT 107.660 533.120 111.200 534.240 ;
  LAYER ME2 ;
  RECT 107.660 533.120 111.200 534.240 ;
  LAYER ME1 ;
  RECT 107.660 533.120 111.200 534.240 ;
 END
 PORT
  LAYER ME4 ;
  RECT 98.980 533.120 102.520 534.240 ;
  LAYER ME3 ;
  RECT 98.980 533.120 102.520 534.240 ;
  LAYER ME2 ;
  RECT 98.980 533.120 102.520 534.240 ;
  LAYER ME1 ;
  RECT 98.980 533.120 102.520 534.240 ;
 END
 PORT
  LAYER ME4 ;
  RECT 55.580 533.120 59.120 534.240 ;
  LAYER ME3 ;
  RECT 55.580 533.120 59.120 534.240 ;
  LAYER ME2 ;
  RECT 55.580 533.120 59.120 534.240 ;
  LAYER ME1 ;
  RECT 55.580 533.120 59.120 534.240 ;
 END
 PORT
  LAYER ME4 ;
  RECT 46.900 533.120 50.440 534.240 ;
  LAYER ME3 ;
  RECT 46.900 533.120 50.440 534.240 ;
  LAYER ME2 ;
  RECT 46.900 533.120 50.440 534.240 ;
  LAYER ME1 ;
  RECT 46.900 533.120 50.440 534.240 ;
 END
 PORT
  LAYER ME4 ;
  RECT 38.220 533.120 41.760 534.240 ;
  LAYER ME3 ;
  RECT 38.220 533.120 41.760 534.240 ;
  LAYER ME2 ;
  RECT 38.220 533.120 41.760 534.240 ;
  LAYER ME1 ;
  RECT 38.220 533.120 41.760 534.240 ;
 END
 PORT
  LAYER ME4 ;
  RECT 29.540 533.120 33.080 534.240 ;
  LAYER ME3 ;
  RECT 29.540 533.120 33.080 534.240 ;
  LAYER ME2 ;
  RECT 29.540 533.120 33.080 534.240 ;
  LAYER ME1 ;
  RECT 29.540 533.120 33.080 534.240 ;
 END
 PORT
  LAYER ME4 ;
  RECT 20.860 533.120 24.400 534.240 ;
  LAYER ME3 ;
  RECT 20.860 533.120 24.400 534.240 ;
  LAYER ME2 ;
  RECT 20.860 533.120 24.400 534.240 ;
  LAYER ME1 ;
  RECT 20.860 533.120 24.400 534.240 ;
 END
 PORT
  LAYER ME4 ;
  RECT 12.180 533.120 15.720 534.240 ;
  LAYER ME3 ;
  RECT 12.180 533.120 15.720 534.240 ;
  LAYER ME2 ;
  RECT 12.180 533.120 15.720 534.240 ;
  LAYER ME1 ;
  RECT 12.180 533.120 15.720 534.240 ;
 END
 PORT
  LAYER ME4 ;
  RECT 334.580 0.000 338.120 1.120 ;
  LAYER ME3 ;
  RECT 334.580 0.000 338.120 1.120 ;
  LAYER ME2 ;
  RECT 334.580 0.000 338.120 1.120 ;
  LAYER ME1 ;
  RECT 334.580 0.000 338.120 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 317.840 0.000 321.380 1.120 ;
  LAYER ME3 ;
  RECT 317.840 0.000 321.380 1.120 ;
  LAYER ME2 ;
  RECT 317.840 0.000 321.380 1.120 ;
  LAYER ME1 ;
  RECT 317.840 0.000 321.380 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 291.180 0.000 294.720 1.120 ;
  LAYER ME3 ;
  RECT 291.180 0.000 294.720 1.120 ;
  LAYER ME2 ;
  RECT 291.180 0.000 294.720 1.120 ;
  LAYER ME1 ;
  RECT 291.180 0.000 294.720 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 269.480 0.000 273.020 1.120 ;
  LAYER ME3 ;
  RECT 269.480 0.000 273.020 1.120 ;
  LAYER ME2 ;
  RECT 269.480 0.000 273.020 1.120 ;
  LAYER ME1 ;
  RECT 269.480 0.000 273.020 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 247.780 0.000 251.320 1.120 ;
  LAYER ME3 ;
  RECT 247.780 0.000 251.320 1.120 ;
  LAYER ME2 ;
  RECT 247.780 0.000 251.320 1.120 ;
  LAYER ME1 ;
  RECT 247.780 0.000 251.320 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 221.120 0.000 224.660 1.120 ;
  LAYER ME3 ;
  RECT 221.120 0.000 224.660 1.120 ;
  LAYER ME2 ;
  RECT 221.120 0.000 224.660 1.120 ;
  LAYER ME1 ;
  RECT 221.120 0.000 224.660 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 135.560 0.000 139.100 1.120 ;
  LAYER ME3 ;
  RECT 135.560 0.000 139.100 1.120 ;
  LAYER ME2 ;
  RECT 135.560 0.000 139.100 1.120 ;
  LAYER ME1 ;
  RECT 135.560 0.000 139.100 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 113.860 0.000 117.400 1.120 ;
  LAYER ME3 ;
  RECT 113.860 0.000 117.400 1.120 ;
  LAYER ME2 ;
  RECT 113.860 0.000 117.400 1.120 ;
  LAYER ME1 ;
  RECT 113.860 0.000 117.400 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 92.160 0.000 95.700 1.120 ;
  LAYER ME3 ;
  RECT 92.160 0.000 95.700 1.120 ;
  LAYER ME2 ;
  RECT 92.160 0.000 95.700 1.120 ;
  LAYER ME1 ;
  RECT 92.160 0.000 95.700 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 70.460 0.000 74.000 1.120 ;
  LAYER ME3 ;
  RECT 70.460 0.000 74.000 1.120 ;
  LAYER ME2 ;
  RECT 70.460 0.000 74.000 1.120 ;
  LAYER ME1 ;
  RECT 70.460 0.000 74.000 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 43.800 0.000 47.340 1.120 ;
  LAYER ME3 ;
  RECT 43.800 0.000 47.340 1.120 ;
  LAYER ME2 ;
  RECT 43.800 0.000 47.340 1.120 ;
  LAYER ME1 ;
  RECT 43.800 0.000 47.340 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 27.060 0.000 30.600 1.120 ;
  LAYER ME3 ;
  RECT 27.060 0.000 30.600 1.120 ;
  LAYER ME2 ;
  RECT 27.060 0.000 30.600 1.120 ;
  LAYER ME1 ;
  RECT 27.060 0.000 30.600 1.120 ;
 END
END GND
PIN VCC
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
 PORT
  LAYER ME4 ;
  RECT 396.300 517.780 397.420 521.020 ;
  LAYER ME3 ;
  RECT 396.300 517.780 397.420 521.020 ;
  LAYER ME2 ;
  RECT 396.300 517.780 397.420 521.020 ;
  LAYER ME1 ;
  RECT 396.300 517.780 397.420 521.020 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 509.940 397.420 513.180 ;
  LAYER ME3 ;
  RECT 396.300 509.940 397.420 513.180 ;
  LAYER ME2 ;
  RECT 396.300 509.940 397.420 513.180 ;
  LAYER ME1 ;
  RECT 396.300 509.940 397.420 513.180 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 502.100 397.420 505.340 ;
  LAYER ME3 ;
  RECT 396.300 502.100 397.420 505.340 ;
  LAYER ME2 ;
  RECT 396.300 502.100 397.420 505.340 ;
  LAYER ME1 ;
  RECT 396.300 502.100 397.420 505.340 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 494.260 397.420 497.500 ;
  LAYER ME3 ;
  RECT 396.300 494.260 397.420 497.500 ;
  LAYER ME2 ;
  RECT 396.300 494.260 397.420 497.500 ;
  LAYER ME1 ;
  RECT 396.300 494.260 397.420 497.500 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 486.420 397.420 489.660 ;
  LAYER ME3 ;
  RECT 396.300 486.420 397.420 489.660 ;
  LAYER ME2 ;
  RECT 396.300 486.420 397.420 489.660 ;
  LAYER ME1 ;
  RECT 396.300 486.420 397.420 489.660 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 478.580 397.420 481.820 ;
  LAYER ME3 ;
  RECT 396.300 478.580 397.420 481.820 ;
  LAYER ME2 ;
  RECT 396.300 478.580 397.420 481.820 ;
  LAYER ME1 ;
  RECT 396.300 478.580 397.420 481.820 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 439.380 397.420 442.620 ;
  LAYER ME3 ;
  RECT 396.300 439.380 397.420 442.620 ;
  LAYER ME2 ;
  RECT 396.300 439.380 397.420 442.620 ;
  LAYER ME1 ;
  RECT 396.300 439.380 397.420 442.620 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 431.540 397.420 434.780 ;
  LAYER ME3 ;
  RECT 396.300 431.540 397.420 434.780 ;
  LAYER ME2 ;
  RECT 396.300 431.540 397.420 434.780 ;
  LAYER ME1 ;
  RECT 396.300 431.540 397.420 434.780 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 423.700 397.420 426.940 ;
  LAYER ME3 ;
  RECT 396.300 423.700 397.420 426.940 ;
  LAYER ME2 ;
  RECT 396.300 423.700 397.420 426.940 ;
  LAYER ME1 ;
  RECT 396.300 423.700 397.420 426.940 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 415.860 397.420 419.100 ;
  LAYER ME3 ;
  RECT 396.300 415.860 397.420 419.100 ;
  LAYER ME2 ;
  RECT 396.300 415.860 397.420 419.100 ;
  LAYER ME1 ;
  RECT 396.300 415.860 397.420 419.100 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 408.020 397.420 411.260 ;
  LAYER ME3 ;
  RECT 396.300 408.020 397.420 411.260 ;
  LAYER ME2 ;
  RECT 396.300 408.020 397.420 411.260 ;
  LAYER ME1 ;
  RECT 396.300 408.020 397.420 411.260 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 400.180 397.420 403.420 ;
  LAYER ME3 ;
  RECT 396.300 400.180 397.420 403.420 ;
  LAYER ME2 ;
  RECT 396.300 400.180 397.420 403.420 ;
  LAYER ME1 ;
  RECT 396.300 400.180 397.420 403.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 360.980 397.420 364.220 ;
  LAYER ME3 ;
  RECT 396.300 360.980 397.420 364.220 ;
  LAYER ME2 ;
  RECT 396.300 360.980 397.420 364.220 ;
  LAYER ME1 ;
  RECT 396.300 360.980 397.420 364.220 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 353.140 397.420 356.380 ;
  LAYER ME3 ;
  RECT 396.300 353.140 397.420 356.380 ;
  LAYER ME2 ;
  RECT 396.300 353.140 397.420 356.380 ;
  LAYER ME1 ;
  RECT 396.300 353.140 397.420 356.380 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 345.300 397.420 348.540 ;
  LAYER ME3 ;
  RECT 396.300 345.300 397.420 348.540 ;
  LAYER ME2 ;
  RECT 396.300 345.300 397.420 348.540 ;
  LAYER ME1 ;
  RECT 396.300 345.300 397.420 348.540 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 337.460 397.420 340.700 ;
  LAYER ME3 ;
  RECT 396.300 337.460 397.420 340.700 ;
  LAYER ME2 ;
  RECT 396.300 337.460 397.420 340.700 ;
  LAYER ME1 ;
  RECT 396.300 337.460 397.420 340.700 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 329.620 397.420 332.860 ;
  LAYER ME3 ;
  RECT 396.300 329.620 397.420 332.860 ;
  LAYER ME2 ;
  RECT 396.300 329.620 397.420 332.860 ;
  LAYER ME1 ;
  RECT 396.300 329.620 397.420 332.860 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 321.780 397.420 325.020 ;
  LAYER ME3 ;
  RECT 396.300 321.780 397.420 325.020 ;
  LAYER ME2 ;
  RECT 396.300 321.780 397.420 325.020 ;
  LAYER ME1 ;
  RECT 396.300 321.780 397.420 325.020 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 282.580 397.420 285.820 ;
  LAYER ME3 ;
  RECT 396.300 282.580 397.420 285.820 ;
  LAYER ME2 ;
  RECT 396.300 282.580 397.420 285.820 ;
  LAYER ME1 ;
  RECT 396.300 282.580 397.420 285.820 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 274.740 397.420 277.980 ;
  LAYER ME3 ;
  RECT 396.300 274.740 397.420 277.980 ;
  LAYER ME2 ;
  RECT 396.300 274.740 397.420 277.980 ;
  LAYER ME1 ;
  RECT 396.300 274.740 397.420 277.980 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 266.900 397.420 270.140 ;
  LAYER ME3 ;
  RECT 396.300 266.900 397.420 270.140 ;
  LAYER ME2 ;
  RECT 396.300 266.900 397.420 270.140 ;
  LAYER ME1 ;
  RECT 396.300 266.900 397.420 270.140 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 259.060 397.420 262.300 ;
  LAYER ME3 ;
  RECT 396.300 259.060 397.420 262.300 ;
  LAYER ME2 ;
  RECT 396.300 259.060 397.420 262.300 ;
  LAYER ME1 ;
  RECT 396.300 259.060 397.420 262.300 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 251.220 397.420 254.460 ;
  LAYER ME3 ;
  RECT 396.300 251.220 397.420 254.460 ;
  LAYER ME2 ;
  RECT 396.300 251.220 397.420 254.460 ;
  LAYER ME1 ;
  RECT 396.300 251.220 397.420 254.460 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 243.380 397.420 246.620 ;
  LAYER ME3 ;
  RECT 396.300 243.380 397.420 246.620 ;
  LAYER ME2 ;
  RECT 396.300 243.380 397.420 246.620 ;
  LAYER ME1 ;
  RECT 396.300 243.380 397.420 246.620 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 204.180 397.420 207.420 ;
  LAYER ME3 ;
  RECT 396.300 204.180 397.420 207.420 ;
  LAYER ME2 ;
  RECT 396.300 204.180 397.420 207.420 ;
  LAYER ME1 ;
  RECT 396.300 204.180 397.420 207.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 196.340 397.420 199.580 ;
  LAYER ME3 ;
  RECT 396.300 196.340 397.420 199.580 ;
  LAYER ME2 ;
  RECT 396.300 196.340 397.420 199.580 ;
  LAYER ME1 ;
  RECT 396.300 196.340 397.420 199.580 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 188.500 397.420 191.740 ;
  LAYER ME3 ;
  RECT 396.300 188.500 397.420 191.740 ;
  LAYER ME2 ;
  RECT 396.300 188.500 397.420 191.740 ;
  LAYER ME1 ;
  RECT 396.300 188.500 397.420 191.740 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 180.660 397.420 183.900 ;
  LAYER ME3 ;
  RECT 396.300 180.660 397.420 183.900 ;
  LAYER ME2 ;
  RECT 396.300 180.660 397.420 183.900 ;
  LAYER ME1 ;
  RECT 396.300 180.660 397.420 183.900 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 172.820 397.420 176.060 ;
  LAYER ME3 ;
  RECT 396.300 172.820 397.420 176.060 ;
  LAYER ME2 ;
  RECT 396.300 172.820 397.420 176.060 ;
  LAYER ME1 ;
  RECT 396.300 172.820 397.420 176.060 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 164.980 397.420 168.220 ;
  LAYER ME3 ;
  RECT 396.300 164.980 397.420 168.220 ;
  LAYER ME2 ;
  RECT 396.300 164.980 397.420 168.220 ;
  LAYER ME1 ;
  RECT 396.300 164.980 397.420 168.220 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 125.780 397.420 129.020 ;
  LAYER ME3 ;
  RECT 396.300 125.780 397.420 129.020 ;
  LAYER ME2 ;
  RECT 396.300 125.780 397.420 129.020 ;
  LAYER ME1 ;
  RECT 396.300 125.780 397.420 129.020 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 117.940 397.420 121.180 ;
  LAYER ME3 ;
  RECT 396.300 117.940 397.420 121.180 ;
  LAYER ME2 ;
  RECT 396.300 117.940 397.420 121.180 ;
  LAYER ME1 ;
  RECT 396.300 117.940 397.420 121.180 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 110.100 397.420 113.340 ;
  LAYER ME3 ;
  RECT 396.300 110.100 397.420 113.340 ;
  LAYER ME2 ;
  RECT 396.300 110.100 397.420 113.340 ;
  LAYER ME1 ;
  RECT 396.300 110.100 397.420 113.340 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 102.260 397.420 105.500 ;
  LAYER ME3 ;
  RECT 396.300 102.260 397.420 105.500 ;
  LAYER ME2 ;
  RECT 396.300 102.260 397.420 105.500 ;
  LAYER ME1 ;
  RECT 396.300 102.260 397.420 105.500 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 94.420 397.420 97.660 ;
  LAYER ME3 ;
  RECT 396.300 94.420 397.420 97.660 ;
  LAYER ME2 ;
  RECT 396.300 94.420 397.420 97.660 ;
  LAYER ME1 ;
  RECT 396.300 94.420 397.420 97.660 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 86.580 397.420 89.820 ;
  LAYER ME3 ;
  RECT 396.300 86.580 397.420 89.820 ;
  LAYER ME2 ;
  RECT 396.300 86.580 397.420 89.820 ;
  LAYER ME1 ;
  RECT 396.300 86.580 397.420 89.820 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 47.380 397.420 50.620 ;
  LAYER ME3 ;
  RECT 396.300 47.380 397.420 50.620 ;
  LAYER ME2 ;
  RECT 396.300 47.380 397.420 50.620 ;
  LAYER ME1 ;
  RECT 396.300 47.380 397.420 50.620 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 39.540 397.420 42.780 ;
  LAYER ME3 ;
  RECT 396.300 39.540 397.420 42.780 ;
  LAYER ME2 ;
  RECT 396.300 39.540 397.420 42.780 ;
  LAYER ME1 ;
  RECT 396.300 39.540 397.420 42.780 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 31.700 397.420 34.940 ;
  LAYER ME3 ;
  RECT 396.300 31.700 397.420 34.940 ;
  LAYER ME2 ;
  RECT 396.300 31.700 397.420 34.940 ;
  LAYER ME1 ;
  RECT 396.300 31.700 397.420 34.940 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 23.860 397.420 27.100 ;
  LAYER ME3 ;
  RECT 396.300 23.860 397.420 27.100 ;
  LAYER ME2 ;
  RECT 396.300 23.860 397.420 27.100 ;
  LAYER ME1 ;
  RECT 396.300 23.860 397.420 27.100 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 16.020 397.420 19.260 ;
  LAYER ME3 ;
  RECT 396.300 16.020 397.420 19.260 ;
  LAYER ME2 ;
  RECT 396.300 16.020 397.420 19.260 ;
  LAYER ME1 ;
  RECT 396.300 16.020 397.420 19.260 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.300 8.180 397.420 11.420 ;
  LAYER ME3 ;
  RECT 396.300 8.180 397.420 11.420 ;
  LAYER ME2 ;
  RECT 396.300 8.180 397.420 11.420 ;
  LAYER ME1 ;
  RECT 396.300 8.180 397.420 11.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 517.780 1.120 521.020 ;
  LAYER ME3 ;
  RECT 0.000 517.780 1.120 521.020 ;
  LAYER ME2 ;
  RECT 0.000 517.780 1.120 521.020 ;
  LAYER ME1 ;
  RECT 0.000 517.780 1.120 521.020 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 509.940 1.120 513.180 ;
  LAYER ME3 ;
  RECT 0.000 509.940 1.120 513.180 ;
  LAYER ME2 ;
  RECT 0.000 509.940 1.120 513.180 ;
  LAYER ME1 ;
  RECT 0.000 509.940 1.120 513.180 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 502.100 1.120 505.340 ;
  LAYER ME3 ;
  RECT 0.000 502.100 1.120 505.340 ;
  LAYER ME2 ;
  RECT 0.000 502.100 1.120 505.340 ;
  LAYER ME1 ;
  RECT 0.000 502.100 1.120 505.340 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 494.260 1.120 497.500 ;
  LAYER ME3 ;
  RECT 0.000 494.260 1.120 497.500 ;
  LAYER ME2 ;
  RECT 0.000 494.260 1.120 497.500 ;
  LAYER ME1 ;
  RECT 0.000 494.260 1.120 497.500 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 486.420 1.120 489.660 ;
  LAYER ME3 ;
  RECT 0.000 486.420 1.120 489.660 ;
  LAYER ME2 ;
  RECT 0.000 486.420 1.120 489.660 ;
  LAYER ME1 ;
  RECT 0.000 486.420 1.120 489.660 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 478.580 1.120 481.820 ;
  LAYER ME3 ;
  RECT 0.000 478.580 1.120 481.820 ;
  LAYER ME2 ;
  RECT 0.000 478.580 1.120 481.820 ;
  LAYER ME1 ;
  RECT 0.000 478.580 1.120 481.820 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 439.380 1.120 442.620 ;
  LAYER ME3 ;
  RECT 0.000 439.380 1.120 442.620 ;
  LAYER ME2 ;
  RECT 0.000 439.380 1.120 442.620 ;
  LAYER ME1 ;
  RECT 0.000 439.380 1.120 442.620 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 431.540 1.120 434.780 ;
  LAYER ME3 ;
  RECT 0.000 431.540 1.120 434.780 ;
  LAYER ME2 ;
  RECT 0.000 431.540 1.120 434.780 ;
  LAYER ME1 ;
  RECT 0.000 431.540 1.120 434.780 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 423.700 1.120 426.940 ;
  LAYER ME3 ;
  RECT 0.000 423.700 1.120 426.940 ;
  LAYER ME2 ;
  RECT 0.000 423.700 1.120 426.940 ;
  LAYER ME1 ;
  RECT 0.000 423.700 1.120 426.940 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 415.860 1.120 419.100 ;
  LAYER ME3 ;
  RECT 0.000 415.860 1.120 419.100 ;
  LAYER ME2 ;
  RECT 0.000 415.860 1.120 419.100 ;
  LAYER ME1 ;
  RECT 0.000 415.860 1.120 419.100 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 408.020 1.120 411.260 ;
  LAYER ME3 ;
  RECT 0.000 408.020 1.120 411.260 ;
  LAYER ME2 ;
  RECT 0.000 408.020 1.120 411.260 ;
  LAYER ME1 ;
  RECT 0.000 408.020 1.120 411.260 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 400.180 1.120 403.420 ;
  LAYER ME3 ;
  RECT 0.000 400.180 1.120 403.420 ;
  LAYER ME2 ;
  RECT 0.000 400.180 1.120 403.420 ;
  LAYER ME1 ;
  RECT 0.000 400.180 1.120 403.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 360.980 1.120 364.220 ;
  LAYER ME3 ;
  RECT 0.000 360.980 1.120 364.220 ;
  LAYER ME2 ;
  RECT 0.000 360.980 1.120 364.220 ;
  LAYER ME1 ;
  RECT 0.000 360.980 1.120 364.220 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 353.140 1.120 356.380 ;
  LAYER ME3 ;
  RECT 0.000 353.140 1.120 356.380 ;
  LAYER ME2 ;
  RECT 0.000 353.140 1.120 356.380 ;
  LAYER ME1 ;
  RECT 0.000 353.140 1.120 356.380 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 345.300 1.120 348.540 ;
  LAYER ME3 ;
  RECT 0.000 345.300 1.120 348.540 ;
  LAYER ME2 ;
  RECT 0.000 345.300 1.120 348.540 ;
  LAYER ME1 ;
  RECT 0.000 345.300 1.120 348.540 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 337.460 1.120 340.700 ;
  LAYER ME3 ;
  RECT 0.000 337.460 1.120 340.700 ;
  LAYER ME2 ;
  RECT 0.000 337.460 1.120 340.700 ;
  LAYER ME1 ;
  RECT 0.000 337.460 1.120 340.700 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 329.620 1.120 332.860 ;
  LAYER ME3 ;
  RECT 0.000 329.620 1.120 332.860 ;
  LAYER ME2 ;
  RECT 0.000 329.620 1.120 332.860 ;
  LAYER ME1 ;
  RECT 0.000 329.620 1.120 332.860 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 321.780 1.120 325.020 ;
  LAYER ME3 ;
  RECT 0.000 321.780 1.120 325.020 ;
  LAYER ME2 ;
  RECT 0.000 321.780 1.120 325.020 ;
  LAYER ME1 ;
  RECT 0.000 321.780 1.120 325.020 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 282.580 1.120 285.820 ;
  LAYER ME3 ;
  RECT 0.000 282.580 1.120 285.820 ;
  LAYER ME2 ;
  RECT 0.000 282.580 1.120 285.820 ;
  LAYER ME1 ;
  RECT 0.000 282.580 1.120 285.820 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 274.740 1.120 277.980 ;
  LAYER ME3 ;
  RECT 0.000 274.740 1.120 277.980 ;
  LAYER ME2 ;
  RECT 0.000 274.740 1.120 277.980 ;
  LAYER ME1 ;
  RECT 0.000 274.740 1.120 277.980 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 266.900 1.120 270.140 ;
  LAYER ME3 ;
  RECT 0.000 266.900 1.120 270.140 ;
  LAYER ME2 ;
  RECT 0.000 266.900 1.120 270.140 ;
  LAYER ME1 ;
  RECT 0.000 266.900 1.120 270.140 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 259.060 1.120 262.300 ;
  LAYER ME3 ;
  RECT 0.000 259.060 1.120 262.300 ;
  LAYER ME2 ;
  RECT 0.000 259.060 1.120 262.300 ;
  LAYER ME1 ;
  RECT 0.000 259.060 1.120 262.300 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 251.220 1.120 254.460 ;
  LAYER ME3 ;
  RECT 0.000 251.220 1.120 254.460 ;
  LAYER ME2 ;
  RECT 0.000 251.220 1.120 254.460 ;
  LAYER ME1 ;
  RECT 0.000 251.220 1.120 254.460 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 243.380 1.120 246.620 ;
  LAYER ME3 ;
  RECT 0.000 243.380 1.120 246.620 ;
  LAYER ME2 ;
  RECT 0.000 243.380 1.120 246.620 ;
  LAYER ME1 ;
  RECT 0.000 243.380 1.120 246.620 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 204.180 1.120 207.420 ;
  LAYER ME3 ;
  RECT 0.000 204.180 1.120 207.420 ;
  LAYER ME2 ;
  RECT 0.000 204.180 1.120 207.420 ;
  LAYER ME1 ;
  RECT 0.000 204.180 1.120 207.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 196.340 1.120 199.580 ;
  LAYER ME3 ;
  RECT 0.000 196.340 1.120 199.580 ;
  LAYER ME2 ;
  RECT 0.000 196.340 1.120 199.580 ;
  LAYER ME1 ;
  RECT 0.000 196.340 1.120 199.580 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 188.500 1.120 191.740 ;
  LAYER ME3 ;
  RECT 0.000 188.500 1.120 191.740 ;
  LAYER ME2 ;
  RECT 0.000 188.500 1.120 191.740 ;
  LAYER ME1 ;
  RECT 0.000 188.500 1.120 191.740 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 180.660 1.120 183.900 ;
  LAYER ME3 ;
  RECT 0.000 180.660 1.120 183.900 ;
  LAYER ME2 ;
  RECT 0.000 180.660 1.120 183.900 ;
  LAYER ME1 ;
  RECT 0.000 180.660 1.120 183.900 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 172.820 1.120 176.060 ;
  LAYER ME3 ;
  RECT 0.000 172.820 1.120 176.060 ;
  LAYER ME2 ;
  RECT 0.000 172.820 1.120 176.060 ;
  LAYER ME1 ;
  RECT 0.000 172.820 1.120 176.060 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 164.980 1.120 168.220 ;
  LAYER ME3 ;
  RECT 0.000 164.980 1.120 168.220 ;
  LAYER ME2 ;
  RECT 0.000 164.980 1.120 168.220 ;
  LAYER ME1 ;
  RECT 0.000 164.980 1.120 168.220 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 125.780 1.120 129.020 ;
  LAYER ME3 ;
  RECT 0.000 125.780 1.120 129.020 ;
  LAYER ME2 ;
  RECT 0.000 125.780 1.120 129.020 ;
  LAYER ME1 ;
  RECT 0.000 125.780 1.120 129.020 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 117.940 1.120 121.180 ;
  LAYER ME3 ;
  RECT 0.000 117.940 1.120 121.180 ;
  LAYER ME2 ;
  RECT 0.000 117.940 1.120 121.180 ;
  LAYER ME1 ;
  RECT 0.000 117.940 1.120 121.180 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 110.100 1.120 113.340 ;
  LAYER ME3 ;
  RECT 0.000 110.100 1.120 113.340 ;
  LAYER ME2 ;
  RECT 0.000 110.100 1.120 113.340 ;
  LAYER ME1 ;
  RECT 0.000 110.100 1.120 113.340 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 102.260 1.120 105.500 ;
  LAYER ME3 ;
  RECT 0.000 102.260 1.120 105.500 ;
  LAYER ME2 ;
  RECT 0.000 102.260 1.120 105.500 ;
  LAYER ME1 ;
  RECT 0.000 102.260 1.120 105.500 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 94.420 1.120 97.660 ;
  LAYER ME3 ;
  RECT 0.000 94.420 1.120 97.660 ;
  LAYER ME2 ;
  RECT 0.000 94.420 1.120 97.660 ;
  LAYER ME1 ;
  RECT 0.000 94.420 1.120 97.660 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 86.580 1.120 89.820 ;
  LAYER ME3 ;
  RECT 0.000 86.580 1.120 89.820 ;
  LAYER ME2 ;
  RECT 0.000 86.580 1.120 89.820 ;
  LAYER ME1 ;
  RECT 0.000 86.580 1.120 89.820 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 47.380 1.120 50.620 ;
  LAYER ME3 ;
  RECT 0.000 47.380 1.120 50.620 ;
  LAYER ME2 ;
  RECT 0.000 47.380 1.120 50.620 ;
  LAYER ME1 ;
  RECT 0.000 47.380 1.120 50.620 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 39.540 1.120 42.780 ;
  LAYER ME3 ;
  RECT 0.000 39.540 1.120 42.780 ;
  LAYER ME2 ;
  RECT 0.000 39.540 1.120 42.780 ;
  LAYER ME1 ;
  RECT 0.000 39.540 1.120 42.780 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 31.700 1.120 34.940 ;
  LAYER ME3 ;
  RECT 0.000 31.700 1.120 34.940 ;
  LAYER ME2 ;
  RECT 0.000 31.700 1.120 34.940 ;
  LAYER ME1 ;
  RECT 0.000 31.700 1.120 34.940 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 23.860 1.120 27.100 ;
  LAYER ME3 ;
  RECT 0.000 23.860 1.120 27.100 ;
  LAYER ME2 ;
  RECT 0.000 23.860 1.120 27.100 ;
  LAYER ME1 ;
  RECT 0.000 23.860 1.120 27.100 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 16.020 1.120 19.260 ;
  LAYER ME3 ;
  RECT 0.000 16.020 1.120 19.260 ;
  LAYER ME2 ;
  RECT 0.000 16.020 1.120 19.260 ;
  LAYER ME1 ;
  RECT 0.000 16.020 1.120 19.260 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 8.180 1.120 11.420 ;
  LAYER ME3 ;
  RECT 0.000 8.180 1.120 11.420 ;
  LAYER ME2 ;
  RECT 0.000 8.180 1.120 11.420 ;
  LAYER ME1 ;
  RECT 0.000 8.180 1.120 11.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 381.080 533.120 384.620 534.240 ;
  LAYER ME3 ;
  RECT 381.080 533.120 384.620 534.240 ;
  LAYER ME2 ;
  RECT 381.080 533.120 384.620 534.240 ;
  LAYER ME1 ;
  RECT 381.080 533.120 384.620 534.240 ;
 END
 PORT
  LAYER ME4 ;
  RECT 372.400 533.120 375.940 534.240 ;
  LAYER ME3 ;
  RECT 372.400 533.120 375.940 534.240 ;
  LAYER ME2 ;
  RECT 372.400 533.120 375.940 534.240 ;
  LAYER ME1 ;
  RECT 372.400 533.120 375.940 534.240 ;
 END
 PORT
  LAYER ME4 ;
  RECT 363.720 533.120 367.260 534.240 ;
  LAYER ME3 ;
  RECT 363.720 533.120 367.260 534.240 ;
  LAYER ME2 ;
  RECT 363.720 533.120 367.260 534.240 ;
  LAYER ME1 ;
  RECT 363.720 533.120 367.260 534.240 ;
 END
 PORT
  LAYER ME4 ;
  RECT 355.040 533.120 358.580 534.240 ;
  LAYER ME3 ;
  RECT 355.040 533.120 358.580 534.240 ;
  LAYER ME2 ;
  RECT 355.040 533.120 358.580 534.240 ;
  LAYER ME1 ;
  RECT 355.040 533.120 358.580 534.240 ;
 END
 PORT
  LAYER ME4 ;
  RECT 311.640 533.120 315.180 534.240 ;
  LAYER ME3 ;
  RECT 311.640 533.120 315.180 534.240 ;
  LAYER ME2 ;
  RECT 311.640 533.120 315.180 534.240 ;
  LAYER ME1 ;
  RECT 311.640 533.120 315.180 534.240 ;
 END
 PORT
  LAYER ME4 ;
  RECT 302.960 533.120 306.500 534.240 ;
  LAYER ME3 ;
  RECT 302.960 533.120 306.500 534.240 ;
  LAYER ME2 ;
  RECT 302.960 533.120 306.500 534.240 ;
  LAYER ME1 ;
  RECT 302.960 533.120 306.500 534.240 ;
 END
 PORT
  LAYER ME4 ;
  RECT 294.280 533.120 297.820 534.240 ;
  LAYER ME3 ;
  RECT 294.280 533.120 297.820 534.240 ;
  LAYER ME2 ;
  RECT 294.280 533.120 297.820 534.240 ;
  LAYER ME1 ;
  RECT 294.280 533.120 297.820 534.240 ;
 END
 PORT
  LAYER ME4 ;
  RECT 285.600 533.120 289.140 534.240 ;
  LAYER ME3 ;
  RECT 285.600 533.120 289.140 534.240 ;
  LAYER ME2 ;
  RECT 285.600 533.120 289.140 534.240 ;
  LAYER ME1 ;
  RECT 285.600 533.120 289.140 534.240 ;
 END
 PORT
  LAYER ME4 ;
  RECT 276.920 533.120 280.460 534.240 ;
  LAYER ME3 ;
  RECT 276.920 533.120 280.460 534.240 ;
  LAYER ME2 ;
  RECT 276.920 533.120 280.460 534.240 ;
  LAYER ME1 ;
  RECT 276.920 533.120 280.460 534.240 ;
 END
 PORT
  LAYER ME4 ;
  RECT 268.240 533.120 271.780 534.240 ;
  LAYER ME3 ;
  RECT 268.240 533.120 271.780 534.240 ;
  LAYER ME2 ;
  RECT 268.240 533.120 271.780 534.240 ;
  LAYER ME1 ;
  RECT 268.240 533.120 271.780 534.240 ;
 END
 PORT
  LAYER ME4 ;
  RECT 224.840 533.120 228.380 534.240 ;
  LAYER ME3 ;
  RECT 224.840 533.120 228.380 534.240 ;
  LAYER ME2 ;
  RECT 224.840 533.120 228.380 534.240 ;
  LAYER ME1 ;
  RECT 224.840 533.120 228.380 534.240 ;
 END
 PORT
  LAYER ME4 ;
  RECT 216.160 533.120 219.700 534.240 ;
  LAYER ME3 ;
  RECT 216.160 533.120 219.700 534.240 ;
  LAYER ME2 ;
  RECT 216.160 533.120 219.700 534.240 ;
  LAYER ME1 ;
  RECT 216.160 533.120 219.700 534.240 ;
 END
 PORT
  LAYER ME4 ;
  RECT 207.480 533.120 211.020 534.240 ;
  LAYER ME3 ;
  RECT 207.480 533.120 211.020 534.240 ;
  LAYER ME2 ;
  RECT 207.480 533.120 211.020 534.240 ;
  LAYER ME1 ;
  RECT 207.480 533.120 211.020 534.240 ;
 END
 PORT
  LAYER ME4 ;
  RECT 198.800 533.120 202.340 534.240 ;
  LAYER ME3 ;
  RECT 198.800 533.120 202.340 534.240 ;
  LAYER ME2 ;
  RECT 198.800 533.120 202.340 534.240 ;
  LAYER ME1 ;
  RECT 198.800 533.120 202.340 534.240 ;
 END
 PORT
  LAYER ME4 ;
  RECT 190.120 533.120 193.660 534.240 ;
  LAYER ME3 ;
  RECT 190.120 533.120 193.660 534.240 ;
  LAYER ME2 ;
  RECT 190.120 533.120 193.660 534.240 ;
  LAYER ME1 ;
  RECT 190.120 533.120 193.660 534.240 ;
 END
 PORT
  LAYER ME4 ;
  RECT 181.440 533.120 184.980 534.240 ;
  LAYER ME3 ;
  RECT 181.440 533.120 184.980 534.240 ;
  LAYER ME2 ;
  RECT 181.440 533.120 184.980 534.240 ;
  LAYER ME1 ;
  RECT 181.440 533.120 184.980 534.240 ;
 END
 PORT
  LAYER ME4 ;
  RECT 138.040 533.120 141.580 534.240 ;
  LAYER ME3 ;
  RECT 138.040 533.120 141.580 534.240 ;
  LAYER ME2 ;
  RECT 138.040 533.120 141.580 534.240 ;
  LAYER ME1 ;
  RECT 138.040 533.120 141.580 534.240 ;
 END
 PORT
  LAYER ME4 ;
  RECT 129.360 533.120 132.900 534.240 ;
  LAYER ME3 ;
  RECT 129.360 533.120 132.900 534.240 ;
  LAYER ME2 ;
  RECT 129.360 533.120 132.900 534.240 ;
  LAYER ME1 ;
  RECT 129.360 533.120 132.900 534.240 ;
 END
 PORT
  LAYER ME4 ;
  RECT 120.680 533.120 124.220 534.240 ;
  LAYER ME3 ;
  RECT 120.680 533.120 124.220 534.240 ;
  LAYER ME2 ;
  RECT 120.680 533.120 124.220 534.240 ;
  LAYER ME1 ;
  RECT 120.680 533.120 124.220 534.240 ;
 END
 PORT
  LAYER ME4 ;
  RECT 112.000 533.120 115.540 534.240 ;
  LAYER ME3 ;
  RECT 112.000 533.120 115.540 534.240 ;
  LAYER ME2 ;
  RECT 112.000 533.120 115.540 534.240 ;
  LAYER ME1 ;
  RECT 112.000 533.120 115.540 534.240 ;
 END
 PORT
  LAYER ME4 ;
  RECT 103.320 533.120 106.860 534.240 ;
  LAYER ME3 ;
  RECT 103.320 533.120 106.860 534.240 ;
  LAYER ME2 ;
  RECT 103.320 533.120 106.860 534.240 ;
  LAYER ME1 ;
  RECT 103.320 533.120 106.860 534.240 ;
 END
 PORT
  LAYER ME4 ;
  RECT 94.640 533.120 98.180 534.240 ;
  LAYER ME3 ;
  RECT 94.640 533.120 98.180 534.240 ;
  LAYER ME2 ;
  RECT 94.640 533.120 98.180 534.240 ;
  LAYER ME1 ;
  RECT 94.640 533.120 98.180 534.240 ;
 END
 PORT
  LAYER ME4 ;
  RECT 51.240 533.120 54.780 534.240 ;
  LAYER ME3 ;
  RECT 51.240 533.120 54.780 534.240 ;
  LAYER ME2 ;
  RECT 51.240 533.120 54.780 534.240 ;
  LAYER ME1 ;
  RECT 51.240 533.120 54.780 534.240 ;
 END
 PORT
  LAYER ME4 ;
  RECT 42.560 533.120 46.100 534.240 ;
  LAYER ME3 ;
  RECT 42.560 533.120 46.100 534.240 ;
  LAYER ME2 ;
  RECT 42.560 533.120 46.100 534.240 ;
  LAYER ME1 ;
  RECT 42.560 533.120 46.100 534.240 ;
 END
 PORT
  LAYER ME4 ;
  RECT 33.880 533.120 37.420 534.240 ;
  LAYER ME3 ;
  RECT 33.880 533.120 37.420 534.240 ;
  LAYER ME2 ;
  RECT 33.880 533.120 37.420 534.240 ;
  LAYER ME1 ;
  RECT 33.880 533.120 37.420 534.240 ;
 END
 PORT
  LAYER ME4 ;
  RECT 25.200 533.120 28.740 534.240 ;
  LAYER ME3 ;
  RECT 25.200 533.120 28.740 534.240 ;
  LAYER ME2 ;
  RECT 25.200 533.120 28.740 534.240 ;
  LAYER ME1 ;
  RECT 25.200 533.120 28.740 534.240 ;
 END
 PORT
  LAYER ME4 ;
  RECT 16.520 533.120 20.060 534.240 ;
  LAYER ME3 ;
  RECT 16.520 533.120 20.060 534.240 ;
  LAYER ME2 ;
  RECT 16.520 533.120 20.060 534.240 ;
  LAYER ME1 ;
  RECT 16.520 533.120 20.060 534.240 ;
 END
 PORT
  LAYER ME4 ;
  RECT 7.840 533.120 11.380 534.240 ;
  LAYER ME3 ;
  RECT 7.840 533.120 11.380 534.240 ;
  LAYER ME2 ;
  RECT 7.840 533.120 11.380 534.240 ;
  LAYER ME1 ;
  RECT 7.840 533.120 11.380 534.240 ;
 END
 PORT
  LAYER ME4 ;
  RECT 325.900 0.000 329.440 1.120 ;
  LAYER ME3 ;
  RECT 325.900 0.000 329.440 1.120 ;
  LAYER ME2 ;
  RECT 325.900 0.000 329.440 1.120 ;
  LAYER ME1 ;
  RECT 325.900 0.000 329.440 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 304.200 0.000 307.740 1.120 ;
  LAYER ME3 ;
  RECT 304.200 0.000 307.740 1.120 ;
  LAYER ME2 ;
  RECT 304.200 0.000 307.740 1.120 ;
  LAYER ME1 ;
  RECT 304.200 0.000 307.740 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 278.160 0.000 281.700 1.120 ;
  LAYER ME3 ;
  RECT 278.160 0.000 281.700 1.120 ;
  LAYER ME2 ;
  RECT 278.160 0.000 281.700 1.120 ;
  LAYER ME1 ;
  RECT 278.160 0.000 281.700 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 261.420 0.000 264.960 1.120 ;
  LAYER ME3 ;
  RECT 261.420 0.000 264.960 1.120 ;
  LAYER ME2 ;
  RECT 261.420 0.000 264.960 1.120 ;
  LAYER ME1 ;
  RECT 261.420 0.000 264.960 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 225.460 0.000 229.000 1.120 ;
  LAYER ME3 ;
  RECT 225.460 0.000 229.000 1.120 ;
  LAYER ME2 ;
  RECT 225.460 0.000 229.000 1.120 ;
  LAYER ME1 ;
  RECT 225.460 0.000 229.000 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 216.780 0.000 220.320 1.120 ;
  LAYER ME3 ;
  RECT 216.780 0.000 220.320 1.120 ;
  LAYER ME2 ;
  RECT 216.780 0.000 220.320 1.120 ;
  LAYER ME1 ;
  RECT 216.780 0.000 220.320 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 126.880 0.000 130.420 1.120 ;
  LAYER ME3 ;
  RECT 126.880 0.000 130.420 1.120 ;
  LAYER ME2 ;
  RECT 126.880 0.000 130.420 1.120 ;
  LAYER ME1 ;
  RECT 126.880 0.000 130.420 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 100.220 0.000 103.760 1.120 ;
  LAYER ME3 ;
  RECT 100.220 0.000 103.760 1.120 ;
  LAYER ME2 ;
  RECT 100.220 0.000 103.760 1.120 ;
  LAYER ME1 ;
  RECT 100.220 0.000 103.760 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 83.480 0.000 87.020 1.120 ;
  LAYER ME3 ;
  RECT 83.480 0.000 87.020 1.120 ;
  LAYER ME2 ;
  RECT 83.480 0.000 87.020 1.120 ;
  LAYER ME1 ;
  RECT 83.480 0.000 87.020 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 56.820 0.000 60.360 1.120 ;
  LAYER ME3 ;
  RECT 56.820 0.000 60.360 1.120 ;
  LAYER ME2 ;
  RECT 56.820 0.000 60.360 1.120 ;
  LAYER ME1 ;
  RECT 56.820 0.000 60.360 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 35.740 0.000 39.280 1.120 ;
  LAYER ME3 ;
  RECT 35.740 0.000 39.280 1.120 ;
  LAYER ME2 ;
  RECT 35.740 0.000 39.280 1.120 ;
  LAYER ME1 ;
  RECT 35.740 0.000 39.280 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 14.040 0.000 17.580 1.120 ;
  LAYER ME3 ;
  RECT 14.040 0.000 17.580 1.120 ;
  LAYER ME2 ;
  RECT 14.040 0.000 17.580 1.120 ;
  LAYER ME1 ;
  RECT 14.040 0.000 17.580 1.120 ;
 END
END VCC
PIN DO19
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 383.840 0.000 384.960 1.120 ;
  LAYER ME3 ;
  RECT 383.840 0.000 384.960 1.120 ;
  LAYER ME2 ;
  RECT 383.840 0.000 384.960 1.120 ;
  LAYER ME1 ;
  RECT 383.840 0.000 384.960 1.120 ;
 END
END DO19
PIN DI19
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 375.160 0.000 376.280 1.120 ;
  LAYER ME3 ;
  RECT 375.160 0.000 376.280 1.120 ;
  LAYER ME2 ;
  RECT 375.160 0.000 376.280 1.120 ;
  LAYER ME1 ;
  RECT 375.160 0.000 376.280 1.120 ;
 END
END DI19
PIN DO18
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 367.100 0.000 368.220 1.120 ;
  LAYER ME3 ;
  RECT 367.100 0.000 368.220 1.120 ;
  LAYER ME2 ;
  RECT 367.100 0.000 368.220 1.120 ;
  LAYER ME1 ;
  RECT 367.100 0.000 368.220 1.120 ;
 END
END DO18
PIN DI18
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 359.040 0.000 360.160 1.120 ;
  LAYER ME3 ;
  RECT 359.040 0.000 360.160 1.120 ;
  LAYER ME2 ;
  RECT 359.040 0.000 360.160 1.120 ;
  LAYER ME1 ;
  RECT 359.040 0.000 360.160 1.120 ;
 END
END DI18
PIN DO17
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 354.080 0.000 355.200 1.120 ;
  LAYER ME3 ;
  RECT 354.080 0.000 355.200 1.120 ;
  LAYER ME2 ;
  RECT 354.080 0.000 355.200 1.120 ;
  LAYER ME1 ;
  RECT 354.080 0.000 355.200 1.120 ;
 END
END DO17
PIN DI17
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 345.400 0.000 346.520 1.120 ;
  LAYER ME3 ;
  RECT 345.400 0.000 346.520 1.120 ;
  LAYER ME2 ;
  RECT 345.400 0.000 346.520 1.120 ;
  LAYER ME1 ;
  RECT 345.400 0.000 346.520 1.120 ;
 END
END DI17
PIN DO16
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 340.440 0.000 341.560 1.120 ;
  LAYER ME3 ;
  RECT 340.440 0.000 341.560 1.120 ;
  LAYER ME2 ;
  RECT 340.440 0.000 341.560 1.120 ;
  LAYER ME1 ;
  RECT 340.440 0.000 341.560 1.120 ;
 END
END DO16
PIN DI16
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 332.380 0.000 333.500 1.120 ;
  LAYER ME3 ;
  RECT 332.380 0.000 333.500 1.120 ;
  LAYER ME2 ;
  RECT 332.380 0.000 333.500 1.120 ;
  LAYER ME1 ;
  RECT 332.380 0.000 333.500 1.120 ;
 END
END DI16
PIN DO15
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 323.700 0.000 324.820 1.120 ;
  LAYER ME3 ;
  RECT 323.700 0.000 324.820 1.120 ;
  LAYER ME2 ;
  RECT 323.700 0.000 324.820 1.120 ;
  LAYER ME1 ;
  RECT 323.700 0.000 324.820 1.120 ;
 END
END DO15
PIN DI15
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 315.640 0.000 316.760 1.120 ;
  LAYER ME3 ;
  RECT 315.640 0.000 316.760 1.120 ;
  LAYER ME2 ;
  RECT 315.640 0.000 316.760 1.120 ;
  LAYER ME1 ;
  RECT 315.640 0.000 316.760 1.120 ;
 END
END DI15
PIN DO14
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 310.680 0.000 311.800 1.120 ;
  LAYER ME3 ;
  RECT 310.680 0.000 311.800 1.120 ;
  LAYER ME2 ;
  RECT 310.680 0.000 311.800 1.120 ;
  LAYER ME1 ;
  RECT 310.680 0.000 311.800 1.120 ;
 END
END DO14
PIN DI14
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 302.000 0.000 303.120 1.120 ;
  LAYER ME3 ;
  RECT 302.000 0.000 303.120 1.120 ;
  LAYER ME2 ;
  RECT 302.000 0.000 303.120 1.120 ;
  LAYER ME1 ;
  RECT 302.000 0.000 303.120 1.120 ;
 END
END DI14
PIN DO13
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 297.660 0.000 298.780 1.120 ;
  LAYER ME3 ;
  RECT 297.660 0.000 298.780 1.120 ;
  LAYER ME2 ;
  RECT 297.660 0.000 298.780 1.120 ;
  LAYER ME1 ;
  RECT 297.660 0.000 298.780 1.120 ;
 END
END DO13
PIN DI13
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 288.980 0.000 290.100 1.120 ;
  LAYER ME3 ;
  RECT 288.980 0.000 290.100 1.120 ;
  LAYER ME2 ;
  RECT 288.980 0.000 290.100 1.120 ;
  LAYER ME1 ;
  RECT 288.980 0.000 290.100 1.120 ;
 END
END DI13
PIN DO12
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 284.020 0.000 285.140 1.120 ;
  LAYER ME3 ;
  RECT 284.020 0.000 285.140 1.120 ;
  LAYER ME2 ;
  RECT 284.020 0.000 285.140 1.120 ;
  LAYER ME1 ;
  RECT 284.020 0.000 285.140 1.120 ;
 END
END DO12
PIN DI12
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 275.960 0.000 277.080 1.120 ;
  LAYER ME3 ;
  RECT 275.960 0.000 277.080 1.120 ;
  LAYER ME2 ;
  RECT 275.960 0.000 277.080 1.120 ;
  LAYER ME1 ;
  RECT 275.960 0.000 277.080 1.120 ;
 END
END DI12
PIN DO11
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 267.280 0.000 268.400 1.120 ;
  LAYER ME3 ;
  RECT 267.280 0.000 268.400 1.120 ;
  LAYER ME2 ;
  RECT 267.280 0.000 268.400 1.120 ;
  LAYER ME1 ;
  RECT 267.280 0.000 268.400 1.120 ;
 END
END DO11
PIN DI11
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 259.220 0.000 260.340 1.120 ;
  LAYER ME3 ;
  RECT 259.220 0.000 260.340 1.120 ;
  LAYER ME2 ;
  RECT 259.220 0.000 260.340 1.120 ;
  LAYER ME1 ;
  RECT 259.220 0.000 260.340 1.120 ;
 END
END DI11
PIN DO10
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 254.260 0.000 255.380 1.120 ;
  LAYER ME3 ;
  RECT 254.260 0.000 255.380 1.120 ;
  LAYER ME2 ;
  RECT 254.260 0.000 255.380 1.120 ;
  LAYER ME1 ;
  RECT 254.260 0.000 255.380 1.120 ;
 END
END DO10
PIN DI10
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 245.580 0.000 246.700 1.120 ;
  LAYER ME3 ;
  RECT 245.580 0.000 246.700 1.120 ;
  LAYER ME2 ;
  RECT 245.580 0.000 246.700 1.120 ;
  LAYER ME1 ;
  RECT 245.580 0.000 246.700 1.120 ;
 END
END DI10
PIN A1
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 240.000 0.000 241.120 1.120 ;
  LAYER ME3 ;
  RECT 240.000 0.000 241.120 1.120 ;
  LAYER ME2 ;
  RECT 240.000 0.000 241.120 1.120 ;
  LAYER ME1 ;
  RECT 240.000 0.000 241.120 1.120 ;
 END
END A1
PIN WEB
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER ME4 ;
  RECT 238.140 0.000 239.260 1.120 ;
  LAYER ME3 ;
  RECT 238.140 0.000 239.260 1.120 ;
  LAYER ME2 ;
  RECT 238.140 0.000 239.260 1.120 ;
  LAYER ME1 ;
  RECT 238.140 0.000 239.260 1.120 ;
 END
END WEB
PIN OE
  DIRECTION INPUT ;
  CAPACITANCE 0.033 ;
 PORT
  LAYER ME4 ;
  RECT 233.180 0.000 234.300 1.120 ;
  LAYER ME3 ;
  RECT 233.180 0.000 234.300 1.120 ;
  LAYER ME2 ;
  RECT 233.180 0.000 234.300 1.120 ;
  LAYER ME1 ;
  RECT 233.180 0.000 234.300 1.120 ;
 END
END OE
PIN CS
  DIRECTION INPUT ;
  CAPACITANCE 0.123 ;
 PORT
  LAYER ME4 ;
  RECT 231.320 0.000 232.440 1.120 ;
  LAYER ME3 ;
  RECT 231.320 0.000 232.440 1.120 ;
  LAYER ME2 ;
  RECT 231.320 0.000 232.440 1.120 ;
  LAYER ME1 ;
  RECT 231.320 0.000 232.440 1.120 ;
 END
END CS
PIN A2
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 210.240 0.000 211.360 1.120 ;
  LAYER ME3 ;
  RECT 210.240 0.000 211.360 1.120 ;
  LAYER ME2 ;
  RECT 210.240 0.000 211.360 1.120 ;
  LAYER ME1 ;
  RECT 210.240 0.000 211.360 1.120 ;
 END
END A2
PIN CK
  DIRECTION INPUT ;
  CAPACITANCE 0.063 ;
 PORT
  LAYER ME4 ;
  RECT 207.140 0.000 208.260 1.120 ;
  LAYER ME3 ;
  RECT 207.140 0.000 208.260 1.120 ;
  LAYER ME2 ;
  RECT 207.140 0.000 208.260 1.120 ;
  LAYER ME1 ;
  RECT 207.140 0.000 208.260 1.120 ;
 END
END CK
PIN A0
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 204.660 0.000 205.780 1.120 ;
  LAYER ME3 ;
  RECT 204.660 0.000 205.780 1.120 ;
  LAYER ME2 ;
  RECT 204.660 0.000 205.780 1.120 ;
  LAYER ME1 ;
  RECT 204.660 0.000 205.780 1.120 ;
 END
END A0
PIN A3
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 200.320 0.000 201.440 1.120 ;
  LAYER ME3 ;
  RECT 200.320 0.000 201.440 1.120 ;
  LAYER ME2 ;
  RECT 200.320 0.000 201.440 1.120 ;
  LAYER ME1 ;
  RECT 200.320 0.000 201.440 1.120 ;
 END
END A3
PIN A4
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 192.880 0.000 194.000 1.120 ;
  LAYER ME3 ;
  RECT 192.880 0.000 194.000 1.120 ;
  LAYER ME2 ;
  RECT 192.880 0.000 194.000 1.120 ;
  LAYER ME1 ;
  RECT 192.880 0.000 194.000 1.120 ;
 END
END A4
PIN A5
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 189.780 0.000 190.900 1.120 ;
  LAYER ME3 ;
  RECT 189.780 0.000 190.900 1.120 ;
  LAYER ME2 ;
  RECT 189.780 0.000 190.900 1.120 ;
  LAYER ME1 ;
  RECT 189.780 0.000 190.900 1.120 ;
 END
END A5
PIN A6
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 182.340 0.000 183.460 1.120 ;
  LAYER ME3 ;
  RECT 182.340 0.000 183.460 1.120 ;
  LAYER ME2 ;
  RECT 182.340 0.000 183.460 1.120 ;
  LAYER ME1 ;
  RECT 182.340 0.000 183.460 1.120 ;
 END
END A6
PIN A7
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 179.240 0.000 180.360 1.120 ;
  LAYER ME3 ;
  RECT 179.240 0.000 180.360 1.120 ;
  LAYER ME2 ;
  RECT 179.240 0.000 180.360 1.120 ;
  LAYER ME1 ;
  RECT 179.240 0.000 180.360 1.120 ;
 END
END A7
PIN A8
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 171.800 0.000 172.920 1.120 ;
  LAYER ME3 ;
  RECT 171.800 0.000 172.920 1.120 ;
  LAYER ME2 ;
  RECT 171.800 0.000 172.920 1.120 ;
  LAYER ME1 ;
  RECT 171.800 0.000 172.920 1.120 ;
 END
END A8
PIN A9
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 168.700 0.000 169.820 1.120 ;
  LAYER ME3 ;
  RECT 168.700 0.000 169.820 1.120 ;
  LAYER ME2 ;
  RECT 168.700 0.000 169.820 1.120 ;
  LAYER ME1 ;
  RECT 168.700 0.000 169.820 1.120 ;
 END
END A9
PIN A10
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 161.260 0.000 162.380 1.120 ;
  LAYER ME3 ;
  RECT 161.260 0.000 162.380 1.120 ;
  LAYER ME2 ;
  RECT 161.260 0.000 162.380 1.120 ;
  LAYER ME1 ;
  RECT 161.260 0.000 162.380 1.120 ;
 END
END A10
PIN DO9
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 150.100 0.000 151.220 1.120 ;
  LAYER ME3 ;
  RECT 150.100 0.000 151.220 1.120 ;
  LAYER ME2 ;
  RECT 150.100 0.000 151.220 1.120 ;
  LAYER ME1 ;
  RECT 150.100 0.000 151.220 1.120 ;
 END
END DO9
PIN DI9
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 141.420 0.000 142.540 1.120 ;
  LAYER ME3 ;
  RECT 141.420 0.000 142.540 1.120 ;
  LAYER ME2 ;
  RECT 141.420 0.000 142.540 1.120 ;
  LAYER ME1 ;
  RECT 141.420 0.000 142.540 1.120 ;
 END
END DI9
PIN DO8
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 133.360 0.000 134.480 1.120 ;
  LAYER ME3 ;
  RECT 133.360 0.000 134.480 1.120 ;
  LAYER ME2 ;
  RECT 133.360 0.000 134.480 1.120 ;
  LAYER ME1 ;
  RECT 133.360 0.000 134.480 1.120 ;
 END
END DO8
PIN DI8
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 124.680 0.000 125.800 1.120 ;
  LAYER ME3 ;
  RECT 124.680 0.000 125.800 1.120 ;
  LAYER ME2 ;
  RECT 124.680 0.000 125.800 1.120 ;
  LAYER ME1 ;
  RECT 124.680 0.000 125.800 1.120 ;
 END
END DI8
PIN DO7
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 119.720 0.000 120.840 1.120 ;
  LAYER ME3 ;
  RECT 119.720 0.000 120.840 1.120 ;
  LAYER ME2 ;
  RECT 119.720 0.000 120.840 1.120 ;
  LAYER ME1 ;
  RECT 119.720 0.000 120.840 1.120 ;
 END
END DO7
PIN DI7
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 111.660 0.000 112.780 1.120 ;
  LAYER ME3 ;
  RECT 111.660 0.000 112.780 1.120 ;
  LAYER ME2 ;
  RECT 111.660 0.000 112.780 1.120 ;
  LAYER ME1 ;
  RECT 111.660 0.000 112.780 1.120 ;
 END
END DI7
PIN DO6
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 106.700 0.000 107.820 1.120 ;
  LAYER ME3 ;
  RECT 106.700 0.000 107.820 1.120 ;
  LAYER ME2 ;
  RECT 106.700 0.000 107.820 1.120 ;
  LAYER ME1 ;
  RECT 106.700 0.000 107.820 1.120 ;
 END
END DO6
PIN DI6
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 98.020 0.000 99.140 1.120 ;
  LAYER ME3 ;
  RECT 98.020 0.000 99.140 1.120 ;
  LAYER ME2 ;
  RECT 98.020 0.000 99.140 1.120 ;
  LAYER ME1 ;
  RECT 98.020 0.000 99.140 1.120 ;
 END
END DI6
PIN DO5
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 89.960 0.000 91.080 1.120 ;
  LAYER ME3 ;
  RECT 89.960 0.000 91.080 1.120 ;
  LAYER ME2 ;
  RECT 89.960 0.000 91.080 1.120 ;
  LAYER ME1 ;
  RECT 89.960 0.000 91.080 1.120 ;
 END
END DO5
PIN DI5
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 81.280 0.000 82.400 1.120 ;
  LAYER ME3 ;
  RECT 81.280 0.000 82.400 1.120 ;
  LAYER ME2 ;
  RECT 81.280 0.000 82.400 1.120 ;
  LAYER ME1 ;
  RECT 81.280 0.000 82.400 1.120 ;
 END
END DI5
PIN DO4
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 76.320 0.000 77.440 1.120 ;
  LAYER ME3 ;
  RECT 76.320 0.000 77.440 1.120 ;
  LAYER ME2 ;
  RECT 76.320 0.000 77.440 1.120 ;
  LAYER ME1 ;
  RECT 76.320 0.000 77.440 1.120 ;
 END
END DO4
PIN DI4
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 68.260 0.000 69.380 1.120 ;
  LAYER ME3 ;
  RECT 68.260 0.000 69.380 1.120 ;
  LAYER ME2 ;
  RECT 68.260 0.000 69.380 1.120 ;
  LAYER ME1 ;
  RECT 68.260 0.000 69.380 1.120 ;
 END
END DI4
PIN DO3
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 63.300 0.000 64.420 1.120 ;
  LAYER ME3 ;
  RECT 63.300 0.000 64.420 1.120 ;
  LAYER ME2 ;
  RECT 63.300 0.000 64.420 1.120 ;
  LAYER ME1 ;
  RECT 63.300 0.000 64.420 1.120 ;
 END
END DO3
PIN DI3
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 54.620 0.000 55.740 1.120 ;
  LAYER ME3 ;
  RECT 54.620 0.000 55.740 1.120 ;
  LAYER ME2 ;
  RECT 54.620 0.000 55.740 1.120 ;
  LAYER ME1 ;
  RECT 54.620 0.000 55.740 1.120 ;
 END
END DI3
PIN DO2
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 50.280 0.000 51.400 1.120 ;
  LAYER ME3 ;
  RECT 50.280 0.000 51.400 1.120 ;
  LAYER ME2 ;
  RECT 50.280 0.000 51.400 1.120 ;
  LAYER ME1 ;
  RECT 50.280 0.000 51.400 1.120 ;
 END
END DO2
PIN DI2
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 41.600 0.000 42.720 1.120 ;
  LAYER ME3 ;
  RECT 41.600 0.000 42.720 1.120 ;
  LAYER ME2 ;
  RECT 41.600 0.000 42.720 1.120 ;
  LAYER ME1 ;
  RECT 41.600 0.000 42.720 1.120 ;
 END
END DI2
PIN DO1
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 33.540 0.000 34.660 1.120 ;
  LAYER ME3 ;
  RECT 33.540 0.000 34.660 1.120 ;
  LAYER ME2 ;
  RECT 33.540 0.000 34.660 1.120 ;
  LAYER ME1 ;
  RECT 33.540 0.000 34.660 1.120 ;
 END
END DO1
PIN DI1
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 24.860 0.000 25.980 1.120 ;
  LAYER ME3 ;
  RECT 24.860 0.000 25.980 1.120 ;
  LAYER ME2 ;
  RECT 24.860 0.000 25.980 1.120 ;
  LAYER ME1 ;
  RECT 24.860 0.000 25.980 1.120 ;
 END
END DI1
PIN DO0
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 19.900 0.000 21.020 1.120 ;
  LAYER ME3 ;
  RECT 19.900 0.000 21.020 1.120 ;
  LAYER ME2 ;
  RECT 19.900 0.000 21.020 1.120 ;
  LAYER ME1 ;
  RECT 19.900 0.000 21.020 1.120 ;
 END
END DO0
PIN DI0
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 11.840 0.000 12.960 1.120 ;
  LAYER ME3 ;
  RECT 11.840 0.000 12.960 1.120 ;
  LAYER ME2 ;
  RECT 11.840 0.000 12.960 1.120 ;
  LAYER ME1 ;
  RECT 11.840 0.000 12.960 1.120 ;
 END
END DI0
OBS
  LAYER ME1 SPACING 0.280 ;
  RECT 0.000 0.140 397.420 534.240 ;
  LAYER ME2 SPACING 0.320 ;
  RECT 0.000 0.140 397.420 534.240 ;
  LAYER ME3 SPACING 0.320 ;
  RECT 0.000 0.140 397.420 534.240 ;
  LAYER ME4 SPACING 0.600 ;
  RECT 0.000 0.140 397.420 534.240 ;
  LAYER VI1 ;
  RECT 0.000 0.140 397.420 534.240 ;
  LAYER VI2 ;
  RECT 0.000 0.140 397.420 534.240 ;
  LAYER VI3 ;
  RECT 0.000 0.140 397.420 534.240 ;
END
END SUMA_1296
END LIBRARY



